//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.10.02
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18
//Device Version: C
//Created Time: Sat Sep 14 13:38:26 2024

module inst_mem (dout, ad);

output [15:0] dout;
input [9:0] ad;

wire [0:0] rom16_inst_0_dout;
wire [1:1] rom16_inst_1_dout;
wire [2:2] rom16_inst_2_dout;
wire [3:3] rom16_inst_3_dout;
wire [4:4] rom16_inst_4_dout;
wire [5:5] rom16_inst_5_dout;
wire [6:6] rom16_inst_6_dout;
wire [7:7] rom16_inst_7_dout;
wire [8:8] rom16_inst_8_dout;
wire [9:9] rom16_inst_9_dout;
wire [10:10] rom16_inst_10_dout;
wire [11:11] rom16_inst_11_dout;
wire [12:12] rom16_inst_12_dout;
wire [13:13] rom16_inst_13_dout;
wire [14:14] rom16_inst_14_dout;
wire [15:15] rom16_inst_15_dout;
wire [0:0] rom16_inst_16_dout;
wire [1:1] rom16_inst_17_dout;
wire [2:2] rom16_inst_18_dout;
wire [3:3] rom16_inst_19_dout;
wire [4:4] rom16_inst_20_dout;
wire [5:5] rom16_inst_21_dout;
wire [6:6] rom16_inst_22_dout;
wire [7:7] rom16_inst_23_dout;
wire [8:8] rom16_inst_24_dout;
wire [9:9] rom16_inst_25_dout;
wire [10:10] rom16_inst_26_dout;
wire [11:11] rom16_inst_27_dout;
wire [12:12] rom16_inst_28_dout;
wire [13:13] rom16_inst_29_dout;
wire [14:14] rom16_inst_30_dout;
wire [15:15] rom16_inst_31_dout;
wire [0:0] rom16_inst_32_dout;
wire [1:1] rom16_inst_33_dout;
wire [2:2] rom16_inst_34_dout;
wire [3:3] rom16_inst_35_dout;
wire [4:4] rom16_inst_36_dout;
wire [5:5] rom16_inst_37_dout;
wire [6:6] rom16_inst_38_dout;
wire [7:7] rom16_inst_39_dout;
wire [8:8] rom16_inst_40_dout;
wire [9:9] rom16_inst_41_dout;
wire [10:10] rom16_inst_42_dout;
wire [11:11] rom16_inst_43_dout;
wire [12:12] rom16_inst_44_dout;
wire [13:13] rom16_inst_45_dout;
wire [14:14] rom16_inst_46_dout;
wire [15:15] rom16_inst_47_dout;
wire [0:0] rom16_inst_48_dout;
wire [1:1] rom16_inst_49_dout;
wire [2:2] rom16_inst_50_dout;
wire [3:3] rom16_inst_51_dout;
wire [4:4] rom16_inst_52_dout;
wire [5:5] rom16_inst_53_dout;
wire [6:6] rom16_inst_54_dout;
wire [7:7] rom16_inst_55_dout;
wire [8:8] rom16_inst_56_dout;
wire [9:9] rom16_inst_57_dout;
wire [10:10] rom16_inst_58_dout;
wire [11:11] rom16_inst_59_dout;
wire [12:12] rom16_inst_60_dout;
wire [13:13] rom16_inst_61_dout;
wire [14:14] rom16_inst_62_dout;
wire [15:15] rom16_inst_63_dout;
wire [0:0] rom16_inst_64_dout;
wire [1:1] rom16_inst_65_dout;
wire [2:2] rom16_inst_66_dout;
wire [3:3] rom16_inst_67_dout;
wire [4:4] rom16_inst_68_dout;
wire [5:5] rom16_inst_69_dout;
wire [6:6] rom16_inst_70_dout;
wire [7:7] rom16_inst_71_dout;
wire [8:8] rom16_inst_72_dout;
wire [9:9] rom16_inst_73_dout;
wire [10:10] rom16_inst_74_dout;
wire [11:11] rom16_inst_75_dout;
wire [12:12] rom16_inst_76_dout;
wire [13:13] rom16_inst_77_dout;
wire [14:14] rom16_inst_78_dout;
wire [15:15] rom16_inst_79_dout;
wire [0:0] rom16_inst_80_dout;
wire [1:1] rom16_inst_81_dout;
wire [2:2] rom16_inst_82_dout;
wire [3:3] rom16_inst_83_dout;
wire [4:4] rom16_inst_84_dout;
wire [5:5] rom16_inst_85_dout;
wire [6:6] rom16_inst_86_dout;
wire [7:7] rom16_inst_87_dout;
wire [8:8] rom16_inst_88_dout;
wire [9:9] rom16_inst_89_dout;
wire [10:10] rom16_inst_90_dout;
wire [11:11] rom16_inst_91_dout;
wire [12:12] rom16_inst_92_dout;
wire [13:13] rom16_inst_93_dout;
wire [14:14] rom16_inst_94_dout;
wire [15:15] rom16_inst_95_dout;
wire [0:0] rom16_inst_96_dout;
wire [1:1] rom16_inst_97_dout;
wire [2:2] rom16_inst_98_dout;
wire [3:3] rom16_inst_99_dout;
wire [4:4] rom16_inst_100_dout;
wire [5:5] rom16_inst_101_dout;
wire [6:6] rom16_inst_102_dout;
wire [7:7] rom16_inst_103_dout;
wire [8:8] rom16_inst_104_dout;
wire [9:9] rom16_inst_105_dout;
wire [10:10] rom16_inst_106_dout;
wire [11:11] rom16_inst_107_dout;
wire [12:12] rom16_inst_108_dout;
wire [13:13] rom16_inst_109_dout;
wire [14:14] rom16_inst_110_dout;
wire [15:15] rom16_inst_111_dout;
wire [0:0] rom16_inst_112_dout;
wire [1:1] rom16_inst_113_dout;
wire [2:2] rom16_inst_114_dout;
wire [3:3] rom16_inst_115_dout;
wire [4:4] rom16_inst_116_dout;
wire [5:5] rom16_inst_117_dout;
wire [6:6] rom16_inst_118_dout;
wire [7:7] rom16_inst_119_dout;
wire [8:8] rom16_inst_120_dout;
wire [9:9] rom16_inst_121_dout;
wire [10:10] rom16_inst_122_dout;
wire [11:11] rom16_inst_123_dout;
wire [12:12] rom16_inst_124_dout;
wire [13:13] rom16_inst_125_dout;
wire [14:14] rom16_inst_126_dout;
wire [15:15] rom16_inst_127_dout;
wire [0:0] rom16_inst_128_dout;
wire [1:1] rom16_inst_129_dout;
wire [2:2] rom16_inst_130_dout;
wire [3:3] rom16_inst_131_dout;
wire [4:4] rom16_inst_132_dout;
wire [5:5] rom16_inst_133_dout;
wire [6:6] rom16_inst_134_dout;
wire [7:7] rom16_inst_135_dout;
wire [8:8] rom16_inst_136_dout;
wire [9:9] rom16_inst_137_dout;
wire [10:10] rom16_inst_138_dout;
wire [11:11] rom16_inst_139_dout;
wire [12:12] rom16_inst_140_dout;
wire [13:13] rom16_inst_141_dout;
wire [14:14] rom16_inst_142_dout;
wire [15:15] rom16_inst_143_dout;
wire [0:0] rom16_inst_144_dout;
wire [1:1] rom16_inst_145_dout;
wire [2:2] rom16_inst_146_dout;
wire [3:3] rom16_inst_147_dout;
wire [4:4] rom16_inst_148_dout;
wire [5:5] rom16_inst_149_dout;
wire [6:6] rom16_inst_150_dout;
wire [7:7] rom16_inst_151_dout;
wire [8:8] rom16_inst_152_dout;
wire [9:9] rom16_inst_153_dout;
wire [10:10] rom16_inst_154_dout;
wire [11:11] rom16_inst_155_dout;
wire [12:12] rom16_inst_156_dout;
wire [13:13] rom16_inst_157_dout;
wire [14:14] rom16_inst_158_dout;
wire [15:15] rom16_inst_159_dout;
wire [0:0] rom16_inst_160_dout;
wire [1:1] rom16_inst_161_dout;
wire [2:2] rom16_inst_162_dout;
wire [3:3] rom16_inst_163_dout;
wire [4:4] rom16_inst_164_dout;
wire [5:5] rom16_inst_165_dout;
wire [6:6] rom16_inst_166_dout;
wire [7:7] rom16_inst_167_dout;
wire [8:8] rom16_inst_168_dout;
wire [9:9] rom16_inst_169_dout;
wire [10:10] rom16_inst_170_dout;
wire [11:11] rom16_inst_171_dout;
wire [12:12] rom16_inst_172_dout;
wire [13:13] rom16_inst_173_dout;
wire [14:14] rom16_inst_174_dout;
wire [15:15] rom16_inst_175_dout;
wire [0:0] rom16_inst_176_dout;
wire [1:1] rom16_inst_177_dout;
wire [2:2] rom16_inst_178_dout;
wire [3:3] rom16_inst_179_dout;
wire [4:4] rom16_inst_180_dout;
wire [5:5] rom16_inst_181_dout;
wire [6:6] rom16_inst_182_dout;
wire [7:7] rom16_inst_183_dout;
wire [8:8] rom16_inst_184_dout;
wire [9:9] rom16_inst_185_dout;
wire [10:10] rom16_inst_186_dout;
wire [11:11] rom16_inst_187_dout;
wire [12:12] rom16_inst_188_dout;
wire [13:13] rom16_inst_189_dout;
wire [14:14] rom16_inst_190_dout;
wire [15:15] rom16_inst_191_dout;
wire [0:0] rom16_inst_192_dout;
wire [1:1] rom16_inst_193_dout;
wire [2:2] rom16_inst_194_dout;
wire [3:3] rom16_inst_195_dout;
wire [4:4] rom16_inst_196_dout;
wire [5:5] rom16_inst_197_dout;
wire [6:6] rom16_inst_198_dout;
wire [7:7] rom16_inst_199_dout;
wire [8:8] rom16_inst_200_dout;
wire [9:9] rom16_inst_201_dout;
wire [10:10] rom16_inst_202_dout;
wire [11:11] rom16_inst_203_dout;
wire [12:12] rom16_inst_204_dout;
wire [13:13] rom16_inst_205_dout;
wire [14:14] rom16_inst_206_dout;
wire [15:15] rom16_inst_207_dout;
wire [0:0] rom16_inst_208_dout;
wire [1:1] rom16_inst_209_dout;
wire [2:2] rom16_inst_210_dout;
wire [3:3] rom16_inst_211_dout;
wire [4:4] rom16_inst_212_dout;
wire [5:5] rom16_inst_213_dout;
wire [6:6] rom16_inst_214_dout;
wire [7:7] rom16_inst_215_dout;
wire [8:8] rom16_inst_216_dout;
wire [9:9] rom16_inst_217_dout;
wire [10:10] rom16_inst_218_dout;
wire [11:11] rom16_inst_219_dout;
wire [12:12] rom16_inst_220_dout;
wire [13:13] rom16_inst_221_dout;
wire [14:14] rom16_inst_222_dout;
wire [15:15] rom16_inst_223_dout;
wire [0:0] rom16_inst_224_dout;
wire [1:1] rom16_inst_225_dout;
wire [2:2] rom16_inst_226_dout;
wire [3:3] rom16_inst_227_dout;
wire [4:4] rom16_inst_228_dout;
wire [5:5] rom16_inst_229_dout;
wire [6:6] rom16_inst_230_dout;
wire [7:7] rom16_inst_231_dout;
wire [8:8] rom16_inst_232_dout;
wire [9:9] rom16_inst_233_dout;
wire [10:10] rom16_inst_234_dout;
wire [11:11] rom16_inst_235_dout;
wire [12:12] rom16_inst_236_dout;
wire [13:13] rom16_inst_237_dout;
wire [14:14] rom16_inst_238_dout;
wire [15:15] rom16_inst_239_dout;
wire [0:0] rom16_inst_240_dout;
wire [1:1] rom16_inst_241_dout;
wire [2:2] rom16_inst_242_dout;
wire [3:3] rom16_inst_243_dout;
wire [4:4] rom16_inst_244_dout;
wire [5:5] rom16_inst_245_dout;
wire [6:6] rom16_inst_246_dout;
wire [7:7] rom16_inst_247_dout;
wire [8:8] rom16_inst_248_dout;
wire [9:9] rom16_inst_249_dout;
wire [10:10] rom16_inst_250_dout;
wire [11:11] rom16_inst_251_dout;
wire [12:12] rom16_inst_252_dout;
wire [13:13] rom16_inst_253_dout;
wire [14:14] rom16_inst_254_dout;
wire [15:15] rom16_inst_255_dout;
wire [0:0] rom16_inst_256_dout;
wire [1:1] rom16_inst_257_dout;
wire [2:2] rom16_inst_258_dout;
wire [3:3] rom16_inst_259_dout;
wire [4:4] rom16_inst_260_dout;
wire [5:5] rom16_inst_261_dout;
wire [6:6] rom16_inst_262_dout;
wire [7:7] rom16_inst_263_dout;
wire [8:8] rom16_inst_264_dout;
wire [9:9] rom16_inst_265_dout;
wire [10:10] rom16_inst_266_dout;
wire [11:11] rom16_inst_267_dout;
wire [12:12] rom16_inst_268_dout;
wire [13:13] rom16_inst_269_dout;
wire [14:14] rom16_inst_270_dout;
wire [15:15] rom16_inst_271_dout;
wire [0:0] rom16_inst_272_dout;
wire [1:1] rom16_inst_273_dout;
wire [2:2] rom16_inst_274_dout;
wire [3:3] rom16_inst_275_dout;
wire [4:4] rom16_inst_276_dout;
wire [5:5] rom16_inst_277_dout;
wire [6:6] rom16_inst_278_dout;
wire [7:7] rom16_inst_279_dout;
wire [8:8] rom16_inst_280_dout;
wire [9:9] rom16_inst_281_dout;
wire [10:10] rom16_inst_282_dout;
wire [11:11] rom16_inst_283_dout;
wire [12:12] rom16_inst_284_dout;
wire [13:13] rom16_inst_285_dout;
wire [14:14] rom16_inst_286_dout;
wire [15:15] rom16_inst_287_dout;
wire [0:0] rom16_inst_288_dout;
wire [1:1] rom16_inst_289_dout;
wire [2:2] rom16_inst_290_dout;
wire [3:3] rom16_inst_291_dout;
wire [4:4] rom16_inst_292_dout;
wire [5:5] rom16_inst_293_dout;
wire [6:6] rom16_inst_294_dout;
wire [7:7] rom16_inst_295_dout;
wire [8:8] rom16_inst_296_dout;
wire [9:9] rom16_inst_297_dout;
wire [10:10] rom16_inst_298_dout;
wire [11:11] rom16_inst_299_dout;
wire [12:12] rom16_inst_300_dout;
wire [13:13] rom16_inst_301_dout;
wire [14:14] rom16_inst_302_dout;
wire [15:15] rom16_inst_303_dout;
wire [0:0] rom16_inst_304_dout;
wire [1:1] rom16_inst_305_dout;
wire [2:2] rom16_inst_306_dout;
wire [3:3] rom16_inst_307_dout;
wire [4:4] rom16_inst_308_dout;
wire [5:5] rom16_inst_309_dout;
wire [6:6] rom16_inst_310_dout;
wire [7:7] rom16_inst_311_dout;
wire [8:8] rom16_inst_312_dout;
wire [9:9] rom16_inst_313_dout;
wire [10:10] rom16_inst_314_dout;
wire [11:11] rom16_inst_315_dout;
wire [12:12] rom16_inst_316_dout;
wire [13:13] rom16_inst_317_dout;
wire [14:14] rom16_inst_318_dout;
wire [15:15] rom16_inst_319_dout;
wire [0:0] rom16_inst_320_dout;
wire [1:1] rom16_inst_321_dout;
wire [2:2] rom16_inst_322_dout;
wire [3:3] rom16_inst_323_dout;
wire [4:4] rom16_inst_324_dout;
wire [5:5] rom16_inst_325_dout;
wire [6:6] rom16_inst_326_dout;
wire [7:7] rom16_inst_327_dout;
wire [8:8] rom16_inst_328_dout;
wire [9:9] rom16_inst_329_dout;
wire [10:10] rom16_inst_330_dout;
wire [11:11] rom16_inst_331_dout;
wire [12:12] rom16_inst_332_dout;
wire [13:13] rom16_inst_333_dout;
wire [14:14] rom16_inst_334_dout;
wire [15:15] rom16_inst_335_dout;
wire [0:0] rom16_inst_336_dout;
wire [1:1] rom16_inst_337_dout;
wire [2:2] rom16_inst_338_dout;
wire [3:3] rom16_inst_339_dout;
wire [4:4] rom16_inst_340_dout;
wire [5:5] rom16_inst_341_dout;
wire [6:6] rom16_inst_342_dout;
wire [7:7] rom16_inst_343_dout;
wire [8:8] rom16_inst_344_dout;
wire [9:9] rom16_inst_345_dout;
wire [10:10] rom16_inst_346_dout;
wire [11:11] rom16_inst_347_dout;
wire [12:12] rom16_inst_348_dout;
wire [13:13] rom16_inst_349_dout;
wire [14:14] rom16_inst_350_dout;
wire [15:15] rom16_inst_351_dout;
wire [0:0] rom16_inst_352_dout;
wire [1:1] rom16_inst_353_dout;
wire [2:2] rom16_inst_354_dout;
wire [3:3] rom16_inst_355_dout;
wire [4:4] rom16_inst_356_dout;
wire [5:5] rom16_inst_357_dout;
wire [6:6] rom16_inst_358_dout;
wire [7:7] rom16_inst_359_dout;
wire [8:8] rom16_inst_360_dout;
wire [9:9] rom16_inst_361_dout;
wire [10:10] rom16_inst_362_dout;
wire [11:11] rom16_inst_363_dout;
wire [12:12] rom16_inst_364_dout;
wire [13:13] rom16_inst_365_dout;
wire [14:14] rom16_inst_366_dout;
wire [15:15] rom16_inst_367_dout;
wire [0:0] rom16_inst_368_dout;
wire [1:1] rom16_inst_369_dout;
wire [2:2] rom16_inst_370_dout;
wire [3:3] rom16_inst_371_dout;
wire [4:4] rom16_inst_372_dout;
wire [5:5] rom16_inst_373_dout;
wire [6:6] rom16_inst_374_dout;
wire [7:7] rom16_inst_375_dout;
wire [8:8] rom16_inst_376_dout;
wire [9:9] rom16_inst_377_dout;
wire [10:10] rom16_inst_378_dout;
wire [11:11] rom16_inst_379_dout;
wire [12:12] rom16_inst_380_dout;
wire [13:13] rom16_inst_381_dout;
wire [14:14] rom16_inst_382_dout;
wire [15:15] rom16_inst_383_dout;
wire [0:0] rom16_inst_384_dout;
wire [1:1] rom16_inst_385_dout;
wire [2:2] rom16_inst_386_dout;
wire [3:3] rom16_inst_387_dout;
wire [4:4] rom16_inst_388_dout;
wire [5:5] rom16_inst_389_dout;
wire [6:6] rom16_inst_390_dout;
wire [7:7] rom16_inst_391_dout;
wire [8:8] rom16_inst_392_dout;
wire [9:9] rom16_inst_393_dout;
wire [10:10] rom16_inst_394_dout;
wire [11:11] rom16_inst_395_dout;
wire [12:12] rom16_inst_396_dout;
wire [13:13] rom16_inst_397_dout;
wire [14:14] rom16_inst_398_dout;
wire [15:15] rom16_inst_399_dout;
wire [0:0] rom16_inst_400_dout;
wire [1:1] rom16_inst_401_dout;
wire [2:2] rom16_inst_402_dout;
wire [3:3] rom16_inst_403_dout;
wire [4:4] rom16_inst_404_dout;
wire [5:5] rom16_inst_405_dout;
wire [6:6] rom16_inst_406_dout;
wire [7:7] rom16_inst_407_dout;
wire [8:8] rom16_inst_408_dout;
wire [9:9] rom16_inst_409_dout;
wire [10:10] rom16_inst_410_dout;
wire [11:11] rom16_inst_411_dout;
wire [12:12] rom16_inst_412_dout;
wire [13:13] rom16_inst_413_dout;
wire [14:14] rom16_inst_414_dout;
wire [15:15] rom16_inst_415_dout;
wire [0:0] rom16_inst_416_dout;
wire [1:1] rom16_inst_417_dout;
wire [2:2] rom16_inst_418_dout;
wire [3:3] rom16_inst_419_dout;
wire [4:4] rom16_inst_420_dout;
wire [5:5] rom16_inst_421_dout;
wire [6:6] rom16_inst_422_dout;
wire [7:7] rom16_inst_423_dout;
wire [8:8] rom16_inst_424_dout;
wire [9:9] rom16_inst_425_dout;
wire [10:10] rom16_inst_426_dout;
wire [11:11] rom16_inst_427_dout;
wire [12:12] rom16_inst_428_dout;
wire [13:13] rom16_inst_429_dout;
wire [14:14] rom16_inst_430_dout;
wire [15:15] rom16_inst_431_dout;
wire [0:0] rom16_inst_432_dout;
wire [1:1] rom16_inst_433_dout;
wire [2:2] rom16_inst_434_dout;
wire [3:3] rom16_inst_435_dout;
wire [4:4] rom16_inst_436_dout;
wire [5:5] rom16_inst_437_dout;
wire [6:6] rom16_inst_438_dout;
wire [7:7] rom16_inst_439_dout;
wire [8:8] rom16_inst_440_dout;
wire [9:9] rom16_inst_441_dout;
wire [10:10] rom16_inst_442_dout;
wire [11:11] rom16_inst_443_dout;
wire [12:12] rom16_inst_444_dout;
wire [13:13] rom16_inst_445_dout;
wire [14:14] rom16_inst_446_dout;
wire [15:15] rom16_inst_447_dout;
wire [0:0] rom16_inst_448_dout;
wire [1:1] rom16_inst_449_dout;
wire [2:2] rom16_inst_450_dout;
wire [3:3] rom16_inst_451_dout;
wire [4:4] rom16_inst_452_dout;
wire [5:5] rom16_inst_453_dout;
wire [6:6] rom16_inst_454_dout;
wire [7:7] rom16_inst_455_dout;
wire [8:8] rom16_inst_456_dout;
wire [9:9] rom16_inst_457_dout;
wire [10:10] rom16_inst_458_dout;
wire [11:11] rom16_inst_459_dout;
wire [12:12] rom16_inst_460_dout;
wire [13:13] rom16_inst_461_dout;
wire [14:14] rom16_inst_462_dout;
wire [15:15] rom16_inst_463_dout;
wire [0:0] rom16_inst_464_dout;
wire [1:1] rom16_inst_465_dout;
wire [2:2] rom16_inst_466_dout;
wire [3:3] rom16_inst_467_dout;
wire [4:4] rom16_inst_468_dout;
wire [5:5] rom16_inst_469_dout;
wire [6:6] rom16_inst_470_dout;
wire [7:7] rom16_inst_471_dout;
wire [8:8] rom16_inst_472_dout;
wire [9:9] rom16_inst_473_dout;
wire [10:10] rom16_inst_474_dout;
wire [11:11] rom16_inst_475_dout;
wire [12:12] rom16_inst_476_dout;
wire [13:13] rom16_inst_477_dout;
wire [14:14] rom16_inst_478_dout;
wire [15:15] rom16_inst_479_dout;
wire [0:0] rom16_inst_480_dout;
wire [1:1] rom16_inst_481_dout;
wire [2:2] rom16_inst_482_dout;
wire [3:3] rom16_inst_483_dout;
wire [4:4] rom16_inst_484_dout;
wire [5:5] rom16_inst_485_dout;
wire [6:6] rom16_inst_486_dout;
wire [7:7] rom16_inst_487_dout;
wire [8:8] rom16_inst_488_dout;
wire [9:9] rom16_inst_489_dout;
wire [10:10] rom16_inst_490_dout;
wire [11:11] rom16_inst_491_dout;
wire [12:12] rom16_inst_492_dout;
wire [13:13] rom16_inst_493_dout;
wire [14:14] rom16_inst_494_dout;
wire [15:15] rom16_inst_495_dout;
wire [0:0] rom16_inst_496_dout;
wire [1:1] rom16_inst_497_dout;
wire [2:2] rom16_inst_498_dout;
wire [3:3] rom16_inst_499_dout;
wire [4:4] rom16_inst_500_dout;
wire [5:5] rom16_inst_501_dout;
wire [6:6] rom16_inst_502_dout;
wire [7:7] rom16_inst_503_dout;
wire [8:8] rom16_inst_504_dout;
wire [9:9] rom16_inst_505_dout;
wire [10:10] rom16_inst_506_dout;
wire [11:11] rom16_inst_507_dout;
wire [12:12] rom16_inst_508_dout;
wire [13:13] rom16_inst_509_dout;
wire [14:14] rom16_inst_510_dout;
wire [15:15] rom16_inst_511_dout;
wire [0:0] rom16_inst_512_dout;
wire [1:1] rom16_inst_513_dout;
wire [2:2] rom16_inst_514_dout;
wire [3:3] rom16_inst_515_dout;
wire [4:4] rom16_inst_516_dout;
wire [5:5] rom16_inst_517_dout;
wire [6:6] rom16_inst_518_dout;
wire [7:7] rom16_inst_519_dout;
wire [8:8] rom16_inst_520_dout;
wire [9:9] rom16_inst_521_dout;
wire [10:10] rom16_inst_522_dout;
wire [11:11] rom16_inst_523_dout;
wire [12:12] rom16_inst_524_dout;
wire [13:13] rom16_inst_525_dout;
wire [14:14] rom16_inst_526_dout;
wire [15:15] rom16_inst_527_dout;
wire [0:0] rom16_inst_528_dout;
wire [1:1] rom16_inst_529_dout;
wire [2:2] rom16_inst_530_dout;
wire [3:3] rom16_inst_531_dout;
wire [4:4] rom16_inst_532_dout;
wire [5:5] rom16_inst_533_dout;
wire [6:6] rom16_inst_534_dout;
wire [7:7] rom16_inst_535_dout;
wire [8:8] rom16_inst_536_dout;
wire [9:9] rom16_inst_537_dout;
wire [10:10] rom16_inst_538_dout;
wire [11:11] rom16_inst_539_dout;
wire [12:12] rom16_inst_540_dout;
wire [13:13] rom16_inst_541_dout;
wire [14:14] rom16_inst_542_dout;
wire [15:15] rom16_inst_543_dout;
wire [0:0] rom16_inst_544_dout;
wire [1:1] rom16_inst_545_dout;
wire [2:2] rom16_inst_546_dout;
wire [3:3] rom16_inst_547_dout;
wire [4:4] rom16_inst_548_dout;
wire [5:5] rom16_inst_549_dout;
wire [6:6] rom16_inst_550_dout;
wire [7:7] rom16_inst_551_dout;
wire [8:8] rom16_inst_552_dout;
wire [9:9] rom16_inst_553_dout;
wire [10:10] rom16_inst_554_dout;
wire [11:11] rom16_inst_555_dout;
wire [12:12] rom16_inst_556_dout;
wire [13:13] rom16_inst_557_dout;
wire [14:14] rom16_inst_558_dout;
wire [15:15] rom16_inst_559_dout;
wire [0:0] rom16_inst_560_dout;
wire [1:1] rom16_inst_561_dout;
wire [2:2] rom16_inst_562_dout;
wire [3:3] rom16_inst_563_dout;
wire [4:4] rom16_inst_564_dout;
wire [5:5] rom16_inst_565_dout;
wire [6:6] rom16_inst_566_dout;
wire [7:7] rom16_inst_567_dout;
wire [8:8] rom16_inst_568_dout;
wire [9:9] rom16_inst_569_dout;
wire [10:10] rom16_inst_570_dout;
wire [11:11] rom16_inst_571_dout;
wire [12:12] rom16_inst_572_dout;
wire [13:13] rom16_inst_573_dout;
wire [14:14] rom16_inst_574_dout;
wire [15:15] rom16_inst_575_dout;
wire [0:0] rom16_inst_576_dout;
wire [1:1] rom16_inst_577_dout;
wire [2:2] rom16_inst_578_dout;
wire [3:3] rom16_inst_579_dout;
wire [4:4] rom16_inst_580_dout;
wire [5:5] rom16_inst_581_dout;
wire [6:6] rom16_inst_582_dout;
wire [7:7] rom16_inst_583_dout;
wire [8:8] rom16_inst_584_dout;
wire [9:9] rom16_inst_585_dout;
wire [10:10] rom16_inst_586_dout;
wire [11:11] rom16_inst_587_dout;
wire [12:12] rom16_inst_588_dout;
wire [13:13] rom16_inst_589_dout;
wire [14:14] rom16_inst_590_dout;
wire [15:15] rom16_inst_591_dout;
wire [0:0] rom16_inst_592_dout;
wire [1:1] rom16_inst_593_dout;
wire [2:2] rom16_inst_594_dout;
wire [3:3] rom16_inst_595_dout;
wire [4:4] rom16_inst_596_dout;
wire [5:5] rom16_inst_597_dout;
wire [6:6] rom16_inst_598_dout;
wire [7:7] rom16_inst_599_dout;
wire [8:8] rom16_inst_600_dout;
wire [9:9] rom16_inst_601_dout;
wire [10:10] rom16_inst_602_dout;
wire [11:11] rom16_inst_603_dout;
wire [12:12] rom16_inst_604_dout;
wire [13:13] rom16_inst_605_dout;
wire [14:14] rom16_inst_606_dout;
wire [15:15] rom16_inst_607_dout;
wire [0:0] rom16_inst_608_dout;
wire [1:1] rom16_inst_609_dout;
wire [2:2] rom16_inst_610_dout;
wire [3:3] rom16_inst_611_dout;
wire [4:4] rom16_inst_612_dout;
wire [5:5] rom16_inst_613_dout;
wire [6:6] rom16_inst_614_dout;
wire [7:7] rom16_inst_615_dout;
wire [8:8] rom16_inst_616_dout;
wire [9:9] rom16_inst_617_dout;
wire [10:10] rom16_inst_618_dout;
wire [11:11] rom16_inst_619_dout;
wire [12:12] rom16_inst_620_dout;
wire [13:13] rom16_inst_621_dout;
wire [14:14] rom16_inst_622_dout;
wire [15:15] rom16_inst_623_dout;
wire [0:0] rom16_inst_624_dout;
wire [1:1] rom16_inst_625_dout;
wire [2:2] rom16_inst_626_dout;
wire [3:3] rom16_inst_627_dout;
wire [4:4] rom16_inst_628_dout;
wire [5:5] rom16_inst_629_dout;
wire [6:6] rom16_inst_630_dout;
wire [7:7] rom16_inst_631_dout;
wire [8:8] rom16_inst_632_dout;
wire [9:9] rom16_inst_633_dout;
wire [10:10] rom16_inst_634_dout;
wire [11:11] rom16_inst_635_dout;
wire [12:12] rom16_inst_636_dout;
wire [13:13] rom16_inst_637_dout;
wire [14:14] rom16_inst_638_dout;
wire [15:15] rom16_inst_639_dout;
wire [0:0] rom16_inst_640_dout;
wire [1:1] rom16_inst_641_dout;
wire [2:2] rom16_inst_642_dout;
wire [3:3] rom16_inst_643_dout;
wire [4:4] rom16_inst_644_dout;
wire [5:5] rom16_inst_645_dout;
wire [6:6] rom16_inst_646_dout;
wire [7:7] rom16_inst_647_dout;
wire [8:8] rom16_inst_648_dout;
wire [9:9] rom16_inst_649_dout;
wire [10:10] rom16_inst_650_dout;
wire [11:11] rom16_inst_651_dout;
wire [12:12] rom16_inst_652_dout;
wire [13:13] rom16_inst_653_dout;
wire [14:14] rom16_inst_654_dout;
wire [15:15] rom16_inst_655_dout;
wire [0:0] rom16_inst_656_dout;
wire [1:1] rom16_inst_657_dout;
wire [2:2] rom16_inst_658_dout;
wire [3:3] rom16_inst_659_dout;
wire [4:4] rom16_inst_660_dout;
wire [5:5] rom16_inst_661_dout;
wire [6:6] rom16_inst_662_dout;
wire [7:7] rom16_inst_663_dout;
wire [8:8] rom16_inst_664_dout;
wire [9:9] rom16_inst_665_dout;
wire [10:10] rom16_inst_666_dout;
wire [11:11] rom16_inst_667_dout;
wire [12:12] rom16_inst_668_dout;
wire [13:13] rom16_inst_669_dout;
wire [14:14] rom16_inst_670_dout;
wire [15:15] rom16_inst_671_dout;
wire [0:0] rom16_inst_672_dout;
wire [1:1] rom16_inst_673_dout;
wire [2:2] rom16_inst_674_dout;
wire [3:3] rom16_inst_675_dout;
wire [4:4] rom16_inst_676_dout;
wire [5:5] rom16_inst_677_dout;
wire [6:6] rom16_inst_678_dout;
wire [7:7] rom16_inst_679_dout;
wire [8:8] rom16_inst_680_dout;
wire [9:9] rom16_inst_681_dout;
wire [10:10] rom16_inst_682_dout;
wire [11:11] rom16_inst_683_dout;
wire [12:12] rom16_inst_684_dout;
wire [13:13] rom16_inst_685_dout;
wire [14:14] rom16_inst_686_dout;
wire [15:15] rom16_inst_687_dout;
wire [0:0] rom16_inst_688_dout;
wire [1:1] rom16_inst_689_dout;
wire [2:2] rom16_inst_690_dout;
wire [3:3] rom16_inst_691_dout;
wire [4:4] rom16_inst_692_dout;
wire [5:5] rom16_inst_693_dout;
wire [6:6] rom16_inst_694_dout;
wire [7:7] rom16_inst_695_dout;
wire [8:8] rom16_inst_696_dout;
wire [9:9] rom16_inst_697_dout;
wire [10:10] rom16_inst_698_dout;
wire [11:11] rom16_inst_699_dout;
wire [12:12] rom16_inst_700_dout;
wire [13:13] rom16_inst_701_dout;
wire [14:14] rom16_inst_702_dout;
wire [15:15] rom16_inst_703_dout;
wire [0:0] rom16_inst_704_dout;
wire [1:1] rom16_inst_705_dout;
wire [2:2] rom16_inst_706_dout;
wire [3:3] rom16_inst_707_dout;
wire [4:4] rom16_inst_708_dout;
wire [5:5] rom16_inst_709_dout;
wire [6:6] rom16_inst_710_dout;
wire [7:7] rom16_inst_711_dout;
wire [8:8] rom16_inst_712_dout;
wire [9:9] rom16_inst_713_dout;
wire [10:10] rom16_inst_714_dout;
wire [11:11] rom16_inst_715_dout;
wire [12:12] rom16_inst_716_dout;
wire [13:13] rom16_inst_717_dout;
wire [14:14] rom16_inst_718_dout;
wire [15:15] rom16_inst_719_dout;
wire [0:0] rom16_inst_720_dout;
wire [1:1] rom16_inst_721_dout;
wire [2:2] rom16_inst_722_dout;
wire [3:3] rom16_inst_723_dout;
wire [4:4] rom16_inst_724_dout;
wire [5:5] rom16_inst_725_dout;
wire [6:6] rom16_inst_726_dout;
wire [7:7] rom16_inst_727_dout;
wire [8:8] rom16_inst_728_dout;
wire [9:9] rom16_inst_729_dout;
wire [10:10] rom16_inst_730_dout;
wire [11:11] rom16_inst_731_dout;
wire [12:12] rom16_inst_732_dout;
wire [13:13] rom16_inst_733_dout;
wire [14:14] rom16_inst_734_dout;
wire [15:15] rom16_inst_735_dout;
wire [0:0] rom16_inst_736_dout;
wire [1:1] rom16_inst_737_dout;
wire [2:2] rom16_inst_738_dout;
wire [3:3] rom16_inst_739_dout;
wire [4:4] rom16_inst_740_dout;
wire [5:5] rom16_inst_741_dout;
wire [6:6] rom16_inst_742_dout;
wire [7:7] rom16_inst_743_dout;
wire [8:8] rom16_inst_744_dout;
wire [9:9] rom16_inst_745_dout;
wire [10:10] rom16_inst_746_dout;
wire [11:11] rom16_inst_747_dout;
wire [12:12] rom16_inst_748_dout;
wire [13:13] rom16_inst_749_dout;
wire [14:14] rom16_inst_750_dout;
wire [15:15] rom16_inst_751_dout;
wire [0:0] rom16_inst_752_dout;
wire [1:1] rom16_inst_753_dout;
wire [2:2] rom16_inst_754_dout;
wire [3:3] rom16_inst_755_dout;
wire [4:4] rom16_inst_756_dout;
wire [5:5] rom16_inst_757_dout;
wire [6:6] rom16_inst_758_dout;
wire [7:7] rom16_inst_759_dout;
wire [8:8] rom16_inst_760_dout;
wire [9:9] rom16_inst_761_dout;
wire [10:10] rom16_inst_762_dout;
wire [11:11] rom16_inst_763_dout;
wire [12:12] rom16_inst_764_dout;
wire [13:13] rom16_inst_765_dout;
wire [14:14] rom16_inst_766_dout;
wire [15:15] rom16_inst_767_dout;
wire [0:0] rom16_inst_768_dout;
wire [1:1] rom16_inst_769_dout;
wire [2:2] rom16_inst_770_dout;
wire [3:3] rom16_inst_771_dout;
wire [4:4] rom16_inst_772_dout;
wire [5:5] rom16_inst_773_dout;
wire [6:6] rom16_inst_774_dout;
wire [7:7] rom16_inst_775_dout;
wire [8:8] rom16_inst_776_dout;
wire [9:9] rom16_inst_777_dout;
wire [10:10] rom16_inst_778_dout;
wire [11:11] rom16_inst_779_dout;
wire [12:12] rom16_inst_780_dout;
wire [13:13] rom16_inst_781_dout;
wire [14:14] rom16_inst_782_dout;
wire [15:15] rom16_inst_783_dout;
wire [0:0] rom16_inst_784_dout;
wire [1:1] rom16_inst_785_dout;
wire [2:2] rom16_inst_786_dout;
wire [3:3] rom16_inst_787_dout;
wire [4:4] rom16_inst_788_dout;
wire [5:5] rom16_inst_789_dout;
wire [6:6] rom16_inst_790_dout;
wire [7:7] rom16_inst_791_dout;
wire [8:8] rom16_inst_792_dout;
wire [9:9] rom16_inst_793_dout;
wire [10:10] rom16_inst_794_dout;
wire [11:11] rom16_inst_795_dout;
wire [12:12] rom16_inst_796_dout;
wire [13:13] rom16_inst_797_dout;
wire [14:14] rom16_inst_798_dout;
wire [15:15] rom16_inst_799_dout;
wire [0:0] rom16_inst_800_dout;
wire [1:1] rom16_inst_801_dout;
wire [2:2] rom16_inst_802_dout;
wire [3:3] rom16_inst_803_dout;
wire [4:4] rom16_inst_804_dout;
wire [5:5] rom16_inst_805_dout;
wire [6:6] rom16_inst_806_dout;
wire [7:7] rom16_inst_807_dout;
wire [8:8] rom16_inst_808_dout;
wire [9:9] rom16_inst_809_dout;
wire [10:10] rom16_inst_810_dout;
wire [11:11] rom16_inst_811_dout;
wire [12:12] rom16_inst_812_dout;
wire [13:13] rom16_inst_813_dout;
wire [14:14] rom16_inst_814_dout;
wire [15:15] rom16_inst_815_dout;
wire [0:0] rom16_inst_816_dout;
wire [1:1] rom16_inst_817_dout;
wire [2:2] rom16_inst_818_dout;
wire [3:3] rom16_inst_819_dout;
wire [4:4] rom16_inst_820_dout;
wire [5:5] rom16_inst_821_dout;
wire [6:6] rom16_inst_822_dout;
wire [7:7] rom16_inst_823_dout;
wire [8:8] rom16_inst_824_dout;
wire [9:9] rom16_inst_825_dout;
wire [10:10] rom16_inst_826_dout;
wire [11:11] rom16_inst_827_dout;
wire [12:12] rom16_inst_828_dout;
wire [13:13] rom16_inst_829_dout;
wire [14:14] rom16_inst_830_dout;
wire [15:15] rom16_inst_831_dout;
wire [0:0] rom16_inst_832_dout;
wire [1:1] rom16_inst_833_dout;
wire [2:2] rom16_inst_834_dout;
wire [3:3] rom16_inst_835_dout;
wire [4:4] rom16_inst_836_dout;
wire [5:5] rom16_inst_837_dout;
wire [6:6] rom16_inst_838_dout;
wire [7:7] rom16_inst_839_dout;
wire [8:8] rom16_inst_840_dout;
wire [9:9] rom16_inst_841_dout;
wire [10:10] rom16_inst_842_dout;
wire [11:11] rom16_inst_843_dout;
wire [12:12] rom16_inst_844_dout;
wire [13:13] rom16_inst_845_dout;
wire [14:14] rom16_inst_846_dout;
wire [15:15] rom16_inst_847_dout;
wire [0:0] rom16_inst_848_dout;
wire [1:1] rom16_inst_849_dout;
wire [2:2] rom16_inst_850_dout;
wire [3:3] rom16_inst_851_dout;
wire [4:4] rom16_inst_852_dout;
wire [5:5] rom16_inst_853_dout;
wire [6:6] rom16_inst_854_dout;
wire [7:7] rom16_inst_855_dout;
wire [8:8] rom16_inst_856_dout;
wire [9:9] rom16_inst_857_dout;
wire [10:10] rom16_inst_858_dout;
wire [11:11] rom16_inst_859_dout;
wire [12:12] rom16_inst_860_dout;
wire [13:13] rom16_inst_861_dout;
wire [14:14] rom16_inst_862_dout;
wire [15:15] rom16_inst_863_dout;
wire [0:0] rom16_inst_864_dout;
wire [1:1] rom16_inst_865_dout;
wire [2:2] rom16_inst_866_dout;
wire [3:3] rom16_inst_867_dout;
wire [4:4] rom16_inst_868_dout;
wire [5:5] rom16_inst_869_dout;
wire [6:6] rom16_inst_870_dout;
wire [7:7] rom16_inst_871_dout;
wire [8:8] rom16_inst_872_dout;
wire [9:9] rom16_inst_873_dout;
wire [10:10] rom16_inst_874_dout;
wire [11:11] rom16_inst_875_dout;
wire [12:12] rom16_inst_876_dout;
wire [13:13] rom16_inst_877_dout;
wire [14:14] rom16_inst_878_dout;
wire [15:15] rom16_inst_879_dout;
wire [0:0] rom16_inst_880_dout;
wire [1:1] rom16_inst_881_dout;
wire [2:2] rom16_inst_882_dout;
wire [3:3] rom16_inst_883_dout;
wire [4:4] rom16_inst_884_dout;
wire [5:5] rom16_inst_885_dout;
wire [6:6] rom16_inst_886_dout;
wire [7:7] rom16_inst_887_dout;
wire [8:8] rom16_inst_888_dout;
wire [9:9] rom16_inst_889_dout;
wire [10:10] rom16_inst_890_dout;
wire [11:11] rom16_inst_891_dout;
wire [12:12] rom16_inst_892_dout;
wire [13:13] rom16_inst_893_dout;
wire [14:14] rom16_inst_894_dout;
wire [15:15] rom16_inst_895_dout;
wire [0:0] rom16_inst_896_dout;
wire [1:1] rom16_inst_897_dout;
wire [2:2] rom16_inst_898_dout;
wire [3:3] rom16_inst_899_dout;
wire [4:4] rom16_inst_900_dout;
wire [5:5] rom16_inst_901_dout;
wire [6:6] rom16_inst_902_dout;
wire [7:7] rom16_inst_903_dout;
wire [8:8] rom16_inst_904_dout;
wire [9:9] rom16_inst_905_dout;
wire [10:10] rom16_inst_906_dout;
wire [11:11] rom16_inst_907_dout;
wire [12:12] rom16_inst_908_dout;
wire [13:13] rom16_inst_909_dout;
wire [14:14] rom16_inst_910_dout;
wire [15:15] rom16_inst_911_dout;
wire [0:0] rom16_inst_912_dout;
wire [1:1] rom16_inst_913_dout;
wire [2:2] rom16_inst_914_dout;
wire [3:3] rom16_inst_915_dout;
wire [4:4] rom16_inst_916_dout;
wire [5:5] rom16_inst_917_dout;
wire [6:6] rom16_inst_918_dout;
wire [7:7] rom16_inst_919_dout;
wire [8:8] rom16_inst_920_dout;
wire [9:9] rom16_inst_921_dout;
wire [10:10] rom16_inst_922_dout;
wire [11:11] rom16_inst_923_dout;
wire [12:12] rom16_inst_924_dout;
wire [13:13] rom16_inst_925_dout;
wire [14:14] rom16_inst_926_dout;
wire [15:15] rom16_inst_927_dout;
wire [0:0] rom16_inst_928_dout;
wire [1:1] rom16_inst_929_dout;
wire [2:2] rom16_inst_930_dout;
wire [3:3] rom16_inst_931_dout;
wire [4:4] rom16_inst_932_dout;
wire [5:5] rom16_inst_933_dout;
wire [6:6] rom16_inst_934_dout;
wire [7:7] rom16_inst_935_dout;
wire [8:8] rom16_inst_936_dout;
wire [9:9] rom16_inst_937_dout;
wire [10:10] rom16_inst_938_dout;
wire [11:11] rom16_inst_939_dout;
wire [12:12] rom16_inst_940_dout;
wire [13:13] rom16_inst_941_dout;
wire [14:14] rom16_inst_942_dout;
wire [15:15] rom16_inst_943_dout;
wire [0:0] rom16_inst_944_dout;
wire [1:1] rom16_inst_945_dout;
wire [2:2] rom16_inst_946_dout;
wire [3:3] rom16_inst_947_dout;
wire [4:4] rom16_inst_948_dout;
wire [5:5] rom16_inst_949_dout;
wire [6:6] rom16_inst_950_dout;
wire [7:7] rom16_inst_951_dout;
wire [8:8] rom16_inst_952_dout;
wire [9:9] rom16_inst_953_dout;
wire [10:10] rom16_inst_954_dout;
wire [11:11] rom16_inst_955_dout;
wire [12:12] rom16_inst_956_dout;
wire [13:13] rom16_inst_957_dout;
wire [14:14] rom16_inst_958_dout;
wire [15:15] rom16_inst_959_dout;
wire [0:0] rom16_inst_960_dout;
wire [1:1] rom16_inst_961_dout;
wire [2:2] rom16_inst_962_dout;
wire [3:3] rom16_inst_963_dout;
wire [4:4] rom16_inst_964_dout;
wire [5:5] rom16_inst_965_dout;
wire [6:6] rom16_inst_966_dout;
wire [7:7] rom16_inst_967_dout;
wire [8:8] rom16_inst_968_dout;
wire [9:9] rom16_inst_969_dout;
wire [10:10] rom16_inst_970_dout;
wire [11:11] rom16_inst_971_dout;
wire [12:12] rom16_inst_972_dout;
wire [13:13] rom16_inst_973_dout;
wire [14:14] rom16_inst_974_dout;
wire [15:15] rom16_inst_975_dout;
wire [0:0] rom16_inst_976_dout;
wire [1:1] rom16_inst_977_dout;
wire [2:2] rom16_inst_978_dout;
wire [3:3] rom16_inst_979_dout;
wire [4:4] rom16_inst_980_dout;
wire [5:5] rom16_inst_981_dout;
wire [6:6] rom16_inst_982_dout;
wire [7:7] rom16_inst_983_dout;
wire [8:8] rom16_inst_984_dout;
wire [9:9] rom16_inst_985_dout;
wire [10:10] rom16_inst_986_dout;
wire [11:11] rom16_inst_987_dout;
wire [12:12] rom16_inst_988_dout;
wire [13:13] rom16_inst_989_dout;
wire [14:14] rom16_inst_990_dout;
wire [15:15] rom16_inst_991_dout;
wire [0:0] rom16_inst_992_dout;
wire [1:1] rom16_inst_993_dout;
wire [2:2] rom16_inst_994_dout;
wire [3:3] rom16_inst_995_dout;
wire [4:4] rom16_inst_996_dout;
wire [5:5] rom16_inst_997_dout;
wire [6:6] rom16_inst_998_dout;
wire [7:7] rom16_inst_999_dout;
wire [8:8] rom16_inst_1000_dout;
wire [9:9] rom16_inst_1001_dout;
wire [10:10] rom16_inst_1002_dout;
wire [11:11] rom16_inst_1003_dout;
wire [12:12] rom16_inst_1004_dout;
wire [13:13] rom16_inst_1005_dout;
wire [14:14] rom16_inst_1006_dout;
wire [15:15] rom16_inst_1007_dout;
wire [0:0] rom16_inst_1008_dout;
wire [1:1] rom16_inst_1009_dout;
wire [2:2] rom16_inst_1010_dout;
wire [3:3] rom16_inst_1011_dout;
wire [4:4] rom16_inst_1012_dout;
wire [5:5] rom16_inst_1013_dout;
wire [6:6] rom16_inst_1014_dout;
wire [7:7] rom16_inst_1015_dout;
wire [8:8] rom16_inst_1016_dout;
wire [9:9] rom16_inst_1017_dout;
wire [10:10] rom16_inst_1018_dout;
wire [11:11] rom16_inst_1019_dout;
wire [12:12] rom16_inst_1020_dout;
wire [13:13] rom16_inst_1021_dout;
wire [14:14] rom16_inst_1022_dout;
wire [15:15] rom16_inst_1023_dout;
wire mux_o_0;
wire mux_o_1;
wire mux_o_2;
wire mux_o_3;
wire mux_o_4;
wire mux_o_5;
wire mux_o_6;
wire mux_o_7;
wire mux_o_8;
wire mux_o_9;
wire mux_o_10;
wire mux_o_11;
wire mux_o_12;
wire mux_o_13;
wire mux_o_14;
wire mux_o_15;
wire mux_o_16;
wire mux_o_17;
wire mux_o_18;
wire mux_o_19;
wire mux_o_20;
wire mux_o_21;
wire mux_o_22;
wire mux_o_23;
wire mux_o_24;
wire mux_o_25;
wire mux_o_26;
wire mux_o_27;
wire mux_o_28;
wire mux_o_29;
wire mux_o_30;
wire mux_o_31;
wire mux_o_32;
wire mux_o_33;
wire mux_o_34;
wire mux_o_35;
wire mux_o_36;
wire mux_o_37;
wire mux_o_38;
wire mux_o_39;
wire mux_o_40;
wire mux_o_41;
wire mux_o_42;
wire mux_o_43;
wire mux_o_44;
wire mux_o_45;
wire mux_o_46;
wire mux_o_47;
wire mux_o_48;
wire mux_o_49;
wire mux_o_50;
wire mux_o_51;
wire mux_o_52;
wire mux_o_53;
wire mux_o_54;
wire mux_o_55;
wire mux_o_56;
wire mux_o_57;
wire mux_o_58;
wire mux_o_59;
wire mux_o_60;
wire mux_o_61;
wire mux_o_63;
wire mux_o_64;
wire mux_o_65;
wire mux_o_66;
wire mux_o_67;
wire mux_o_68;
wire mux_o_69;
wire mux_o_70;
wire mux_o_71;
wire mux_o_72;
wire mux_o_73;
wire mux_o_74;
wire mux_o_75;
wire mux_o_76;
wire mux_o_77;
wire mux_o_78;
wire mux_o_79;
wire mux_o_80;
wire mux_o_81;
wire mux_o_82;
wire mux_o_83;
wire mux_o_84;
wire mux_o_85;
wire mux_o_86;
wire mux_o_87;
wire mux_o_88;
wire mux_o_89;
wire mux_o_90;
wire mux_o_91;
wire mux_o_92;
wire mux_o_93;
wire mux_o_94;
wire mux_o_95;
wire mux_o_96;
wire mux_o_97;
wire mux_o_98;
wire mux_o_99;
wire mux_o_100;
wire mux_o_101;
wire mux_o_102;
wire mux_o_103;
wire mux_o_104;
wire mux_o_105;
wire mux_o_106;
wire mux_o_107;
wire mux_o_108;
wire mux_o_109;
wire mux_o_110;
wire mux_o_111;
wire mux_o_112;
wire mux_o_113;
wire mux_o_114;
wire mux_o_115;
wire mux_o_116;
wire mux_o_117;
wire mux_o_118;
wire mux_o_119;
wire mux_o_120;
wire mux_o_121;
wire mux_o_122;
wire mux_o_123;
wire mux_o_124;
wire mux_o_126;
wire mux_o_127;
wire mux_o_128;
wire mux_o_129;
wire mux_o_130;
wire mux_o_131;
wire mux_o_132;
wire mux_o_133;
wire mux_o_134;
wire mux_o_135;
wire mux_o_136;
wire mux_o_137;
wire mux_o_138;
wire mux_o_139;
wire mux_o_140;
wire mux_o_141;
wire mux_o_142;
wire mux_o_143;
wire mux_o_144;
wire mux_o_145;
wire mux_o_146;
wire mux_o_147;
wire mux_o_148;
wire mux_o_149;
wire mux_o_150;
wire mux_o_151;
wire mux_o_152;
wire mux_o_153;
wire mux_o_154;
wire mux_o_155;
wire mux_o_156;
wire mux_o_157;
wire mux_o_158;
wire mux_o_159;
wire mux_o_160;
wire mux_o_161;
wire mux_o_162;
wire mux_o_163;
wire mux_o_164;
wire mux_o_165;
wire mux_o_166;
wire mux_o_167;
wire mux_o_168;
wire mux_o_169;
wire mux_o_170;
wire mux_o_171;
wire mux_o_172;
wire mux_o_173;
wire mux_o_174;
wire mux_o_175;
wire mux_o_176;
wire mux_o_177;
wire mux_o_178;
wire mux_o_179;
wire mux_o_180;
wire mux_o_181;
wire mux_o_182;
wire mux_o_183;
wire mux_o_184;
wire mux_o_185;
wire mux_o_186;
wire mux_o_187;
wire mux_o_189;
wire mux_o_190;
wire mux_o_191;
wire mux_o_192;
wire mux_o_193;
wire mux_o_194;
wire mux_o_195;
wire mux_o_196;
wire mux_o_197;
wire mux_o_198;
wire mux_o_199;
wire mux_o_200;
wire mux_o_201;
wire mux_o_202;
wire mux_o_203;
wire mux_o_204;
wire mux_o_205;
wire mux_o_206;
wire mux_o_207;
wire mux_o_208;
wire mux_o_209;
wire mux_o_210;
wire mux_o_211;
wire mux_o_212;
wire mux_o_213;
wire mux_o_214;
wire mux_o_215;
wire mux_o_216;
wire mux_o_217;
wire mux_o_218;
wire mux_o_219;
wire mux_o_220;
wire mux_o_221;
wire mux_o_222;
wire mux_o_223;
wire mux_o_224;
wire mux_o_225;
wire mux_o_226;
wire mux_o_227;
wire mux_o_228;
wire mux_o_229;
wire mux_o_230;
wire mux_o_231;
wire mux_o_232;
wire mux_o_233;
wire mux_o_234;
wire mux_o_235;
wire mux_o_236;
wire mux_o_237;
wire mux_o_238;
wire mux_o_239;
wire mux_o_240;
wire mux_o_241;
wire mux_o_242;
wire mux_o_243;
wire mux_o_244;
wire mux_o_245;
wire mux_o_246;
wire mux_o_247;
wire mux_o_248;
wire mux_o_249;
wire mux_o_250;
wire mux_o_252;
wire mux_o_253;
wire mux_o_254;
wire mux_o_255;
wire mux_o_256;
wire mux_o_257;
wire mux_o_258;
wire mux_o_259;
wire mux_o_260;
wire mux_o_261;
wire mux_o_262;
wire mux_o_263;
wire mux_o_264;
wire mux_o_265;
wire mux_o_266;
wire mux_o_267;
wire mux_o_268;
wire mux_o_269;
wire mux_o_270;
wire mux_o_271;
wire mux_o_272;
wire mux_o_273;
wire mux_o_274;
wire mux_o_275;
wire mux_o_276;
wire mux_o_277;
wire mux_o_278;
wire mux_o_279;
wire mux_o_280;
wire mux_o_281;
wire mux_o_282;
wire mux_o_283;
wire mux_o_284;
wire mux_o_285;
wire mux_o_286;
wire mux_o_287;
wire mux_o_288;
wire mux_o_289;
wire mux_o_290;
wire mux_o_291;
wire mux_o_292;
wire mux_o_293;
wire mux_o_294;
wire mux_o_295;
wire mux_o_296;
wire mux_o_297;
wire mux_o_298;
wire mux_o_299;
wire mux_o_300;
wire mux_o_301;
wire mux_o_302;
wire mux_o_303;
wire mux_o_304;
wire mux_o_305;
wire mux_o_306;
wire mux_o_307;
wire mux_o_308;
wire mux_o_309;
wire mux_o_310;
wire mux_o_311;
wire mux_o_312;
wire mux_o_313;
wire mux_o_315;
wire mux_o_316;
wire mux_o_317;
wire mux_o_318;
wire mux_o_319;
wire mux_o_320;
wire mux_o_321;
wire mux_o_322;
wire mux_o_323;
wire mux_o_324;
wire mux_o_325;
wire mux_o_326;
wire mux_o_327;
wire mux_o_328;
wire mux_o_329;
wire mux_o_330;
wire mux_o_331;
wire mux_o_332;
wire mux_o_333;
wire mux_o_334;
wire mux_o_335;
wire mux_o_336;
wire mux_o_337;
wire mux_o_338;
wire mux_o_339;
wire mux_o_340;
wire mux_o_341;
wire mux_o_342;
wire mux_o_343;
wire mux_o_344;
wire mux_o_345;
wire mux_o_346;
wire mux_o_347;
wire mux_o_348;
wire mux_o_349;
wire mux_o_350;
wire mux_o_351;
wire mux_o_352;
wire mux_o_353;
wire mux_o_354;
wire mux_o_355;
wire mux_o_356;
wire mux_o_357;
wire mux_o_358;
wire mux_o_359;
wire mux_o_360;
wire mux_o_361;
wire mux_o_362;
wire mux_o_363;
wire mux_o_364;
wire mux_o_365;
wire mux_o_366;
wire mux_o_367;
wire mux_o_368;
wire mux_o_369;
wire mux_o_370;
wire mux_o_371;
wire mux_o_372;
wire mux_o_373;
wire mux_o_374;
wire mux_o_375;
wire mux_o_376;
wire mux_o_378;
wire mux_o_379;
wire mux_o_380;
wire mux_o_381;
wire mux_o_382;
wire mux_o_383;
wire mux_o_384;
wire mux_o_385;
wire mux_o_386;
wire mux_o_387;
wire mux_o_388;
wire mux_o_389;
wire mux_o_390;
wire mux_o_391;
wire mux_o_392;
wire mux_o_393;
wire mux_o_394;
wire mux_o_395;
wire mux_o_396;
wire mux_o_397;
wire mux_o_398;
wire mux_o_399;
wire mux_o_400;
wire mux_o_401;
wire mux_o_402;
wire mux_o_403;
wire mux_o_404;
wire mux_o_405;
wire mux_o_406;
wire mux_o_407;
wire mux_o_408;
wire mux_o_409;
wire mux_o_410;
wire mux_o_411;
wire mux_o_412;
wire mux_o_413;
wire mux_o_414;
wire mux_o_415;
wire mux_o_416;
wire mux_o_417;
wire mux_o_418;
wire mux_o_419;
wire mux_o_420;
wire mux_o_421;
wire mux_o_422;
wire mux_o_423;
wire mux_o_424;
wire mux_o_425;
wire mux_o_426;
wire mux_o_427;
wire mux_o_428;
wire mux_o_429;
wire mux_o_430;
wire mux_o_431;
wire mux_o_432;
wire mux_o_433;
wire mux_o_434;
wire mux_o_435;
wire mux_o_436;
wire mux_o_437;
wire mux_o_438;
wire mux_o_439;
wire mux_o_441;
wire mux_o_442;
wire mux_o_443;
wire mux_o_444;
wire mux_o_445;
wire mux_o_446;
wire mux_o_447;
wire mux_o_448;
wire mux_o_449;
wire mux_o_450;
wire mux_o_451;
wire mux_o_452;
wire mux_o_453;
wire mux_o_454;
wire mux_o_455;
wire mux_o_456;
wire mux_o_457;
wire mux_o_458;
wire mux_o_459;
wire mux_o_460;
wire mux_o_461;
wire mux_o_462;
wire mux_o_463;
wire mux_o_464;
wire mux_o_465;
wire mux_o_466;
wire mux_o_467;
wire mux_o_468;
wire mux_o_469;
wire mux_o_470;
wire mux_o_471;
wire mux_o_472;
wire mux_o_473;
wire mux_o_474;
wire mux_o_475;
wire mux_o_476;
wire mux_o_477;
wire mux_o_478;
wire mux_o_479;
wire mux_o_480;
wire mux_o_481;
wire mux_o_482;
wire mux_o_483;
wire mux_o_484;
wire mux_o_485;
wire mux_o_486;
wire mux_o_487;
wire mux_o_488;
wire mux_o_489;
wire mux_o_490;
wire mux_o_491;
wire mux_o_492;
wire mux_o_493;
wire mux_o_494;
wire mux_o_495;
wire mux_o_496;
wire mux_o_497;
wire mux_o_498;
wire mux_o_499;
wire mux_o_500;
wire mux_o_501;
wire mux_o_502;
wire mux_o_504;
wire mux_o_505;
wire mux_o_506;
wire mux_o_507;
wire mux_o_508;
wire mux_o_509;
wire mux_o_510;
wire mux_o_511;
wire mux_o_512;
wire mux_o_513;
wire mux_o_514;
wire mux_o_515;
wire mux_o_516;
wire mux_o_517;
wire mux_o_518;
wire mux_o_519;
wire mux_o_520;
wire mux_o_521;
wire mux_o_522;
wire mux_o_523;
wire mux_o_524;
wire mux_o_525;
wire mux_o_526;
wire mux_o_527;
wire mux_o_528;
wire mux_o_529;
wire mux_o_530;
wire mux_o_531;
wire mux_o_532;
wire mux_o_533;
wire mux_o_534;
wire mux_o_535;
wire mux_o_536;
wire mux_o_537;
wire mux_o_538;
wire mux_o_539;
wire mux_o_540;
wire mux_o_541;
wire mux_o_542;
wire mux_o_543;
wire mux_o_544;
wire mux_o_545;
wire mux_o_546;
wire mux_o_547;
wire mux_o_548;
wire mux_o_549;
wire mux_o_550;
wire mux_o_551;
wire mux_o_552;
wire mux_o_553;
wire mux_o_554;
wire mux_o_555;
wire mux_o_556;
wire mux_o_557;
wire mux_o_558;
wire mux_o_559;
wire mux_o_560;
wire mux_o_561;
wire mux_o_562;
wire mux_o_563;
wire mux_o_564;
wire mux_o_565;
wire mux_o_567;
wire mux_o_568;
wire mux_o_569;
wire mux_o_570;
wire mux_o_571;
wire mux_o_572;
wire mux_o_573;
wire mux_o_574;
wire mux_o_575;
wire mux_o_576;
wire mux_o_577;
wire mux_o_578;
wire mux_o_579;
wire mux_o_580;
wire mux_o_581;
wire mux_o_582;
wire mux_o_583;
wire mux_o_584;
wire mux_o_585;
wire mux_o_586;
wire mux_o_587;
wire mux_o_588;
wire mux_o_589;
wire mux_o_590;
wire mux_o_591;
wire mux_o_592;
wire mux_o_593;
wire mux_o_594;
wire mux_o_595;
wire mux_o_596;
wire mux_o_597;
wire mux_o_598;
wire mux_o_599;
wire mux_o_600;
wire mux_o_601;
wire mux_o_602;
wire mux_o_603;
wire mux_o_604;
wire mux_o_605;
wire mux_o_606;
wire mux_o_607;
wire mux_o_608;
wire mux_o_609;
wire mux_o_610;
wire mux_o_611;
wire mux_o_612;
wire mux_o_613;
wire mux_o_614;
wire mux_o_615;
wire mux_o_616;
wire mux_o_617;
wire mux_o_618;
wire mux_o_619;
wire mux_o_620;
wire mux_o_621;
wire mux_o_622;
wire mux_o_623;
wire mux_o_624;
wire mux_o_625;
wire mux_o_626;
wire mux_o_627;
wire mux_o_628;
wire mux_o_630;
wire mux_o_631;
wire mux_o_632;
wire mux_o_633;
wire mux_o_634;
wire mux_o_635;
wire mux_o_636;
wire mux_o_637;
wire mux_o_638;
wire mux_o_639;
wire mux_o_640;
wire mux_o_641;
wire mux_o_642;
wire mux_o_643;
wire mux_o_644;
wire mux_o_645;
wire mux_o_646;
wire mux_o_647;
wire mux_o_648;
wire mux_o_649;
wire mux_o_650;
wire mux_o_651;
wire mux_o_652;
wire mux_o_653;
wire mux_o_654;
wire mux_o_655;
wire mux_o_656;
wire mux_o_657;
wire mux_o_658;
wire mux_o_659;
wire mux_o_660;
wire mux_o_661;
wire mux_o_662;
wire mux_o_663;
wire mux_o_664;
wire mux_o_665;
wire mux_o_666;
wire mux_o_667;
wire mux_o_668;
wire mux_o_669;
wire mux_o_670;
wire mux_o_671;
wire mux_o_672;
wire mux_o_673;
wire mux_o_674;
wire mux_o_675;
wire mux_o_676;
wire mux_o_677;
wire mux_o_678;
wire mux_o_679;
wire mux_o_680;
wire mux_o_681;
wire mux_o_682;
wire mux_o_683;
wire mux_o_684;
wire mux_o_685;
wire mux_o_686;
wire mux_o_687;
wire mux_o_688;
wire mux_o_689;
wire mux_o_690;
wire mux_o_691;
wire mux_o_693;
wire mux_o_694;
wire mux_o_695;
wire mux_o_696;
wire mux_o_697;
wire mux_o_698;
wire mux_o_699;
wire mux_o_700;
wire mux_o_701;
wire mux_o_702;
wire mux_o_703;
wire mux_o_704;
wire mux_o_705;
wire mux_o_706;
wire mux_o_707;
wire mux_o_708;
wire mux_o_709;
wire mux_o_710;
wire mux_o_711;
wire mux_o_712;
wire mux_o_713;
wire mux_o_714;
wire mux_o_715;
wire mux_o_716;
wire mux_o_717;
wire mux_o_718;
wire mux_o_719;
wire mux_o_720;
wire mux_o_721;
wire mux_o_722;
wire mux_o_723;
wire mux_o_724;
wire mux_o_725;
wire mux_o_726;
wire mux_o_727;
wire mux_o_728;
wire mux_o_729;
wire mux_o_730;
wire mux_o_731;
wire mux_o_732;
wire mux_o_733;
wire mux_o_734;
wire mux_o_735;
wire mux_o_736;
wire mux_o_737;
wire mux_o_738;
wire mux_o_739;
wire mux_o_740;
wire mux_o_741;
wire mux_o_742;
wire mux_o_743;
wire mux_o_744;
wire mux_o_745;
wire mux_o_746;
wire mux_o_747;
wire mux_o_748;
wire mux_o_749;
wire mux_o_750;
wire mux_o_751;
wire mux_o_752;
wire mux_o_753;
wire mux_o_754;
wire mux_o_756;
wire mux_o_757;
wire mux_o_758;
wire mux_o_759;
wire mux_o_760;
wire mux_o_761;
wire mux_o_762;
wire mux_o_763;
wire mux_o_764;
wire mux_o_765;
wire mux_o_766;
wire mux_o_767;
wire mux_o_768;
wire mux_o_769;
wire mux_o_770;
wire mux_o_771;
wire mux_o_772;
wire mux_o_773;
wire mux_o_774;
wire mux_o_775;
wire mux_o_776;
wire mux_o_777;
wire mux_o_778;
wire mux_o_779;
wire mux_o_780;
wire mux_o_781;
wire mux_o_782;
wire mux_o_783;
wire mux_o_784;
wire mux_o_785;
wire mux_o_786;
wire mux_o_787;
wire mux_o_788;
wire mux_o_789;
wire mux_o_790;
wire mux_o_791;
wire mux_o_792;
wire mux_o_793;
wire mux_o_794;
wire mux_o_795;
wire mux_o_796;
wire mux_o_797;
wire mux_o_798;
wire mux_o_799;
wire mux_o_800;
wire mux_o_801;
wire mux_o_802;
wire mux_o_803;
wire mux_o_804;
wire mux_o_805;
wire mux_o_806;
wire mux_o_807;
wire mux_o_808;
wire mux_o_809;
wire mux_o_810;
wire mux_o_811;
wire mux_o_812;
wire mux_o_813;
wire mux_o_814;
wire mux_o_815;
wire mux_o_816;
wire mux_o_817;
wire mux_o_819;
wire mux_o_820;
wire mux_o_821;
wire mux_o_822;
wire mux_o_823;
wire mux_o_824;
wire mux_o_825;
wire mux_o_826;
wire mux_o_827;
wire mux_o_828;
wire mux_o_829;
wire mux_o_830;
wire mux_o_831;
wire mux_o_832;
wire mux_o_833;
wire mux_o_834;
wire mux_o_835;
wire mux_o_836;
wire mux_o_837;
wire mux_o_838;
wire mux_o_839;
wire mux_o_840;
wire mux_o_841;
wire mux_o_842;
wire mux_o_843;
wire mux_o_844;
wire mux_o_845;
wire mux_o_846;
wire mux_o_847;
wire mux_o_848;
wire mux_o_849;
wire mux_o_850;
wire mux_o_851;
wire mux_o_852;
wire mux_o_853;
wire mux_o_854;
wire mux_o_855;
wire mux_o_856;
wire mux_o_857;
wire mux_o_858;
wire mux_o_859;
wire mux_o_860;
wire mux_o_861;
wire mux_o_862;
wire mux_o_863;
wire mux_o_864;
wire mux_o_865;
wire mux_o_866;
wire mux_o_867;
wire mux_o_868;
wire mux_o_869;
wire mux_o_870;
wire mux_o_871;
wire mux_o_872;
wire mux_o_873;
wire mux_o_874;
wire mux_o_875;
wire mux_o_876;
wire mux_o_877;
wire mux_o_878;
wire mux_o_879;
wire mux_o_880;
wire mux_o_882;
wire mux_o_883;
wire mux_o_884;
wire mux_o_885;
wire mux_o_886;
wire mux_o_887;
wire mux_o_888;
wire mux_o_889;
wire mux_o_890;
wire mux_o_891;
wire mux_o_892;
wire mux_o_893;
wire mux_o_894;
wire mux_o_895;
wire mux_o_896;
wire mux_o_897;
wire mux_o_898;
wire mux_o_899;
wire mux_o_900;
wire mux_o_901;
wire mux_o_902;
wire mux_o_903;
wire mux_o_904;
wire mux_o_905;
wire mux_o_906;
wire mux_o_907;
wire mux_o_908;
wire mux_o_909;
wire mux_o_910;
wire mux_o_911;
wire mux_o_912;
wire mux_o_913;
wire mux_o_914;
wire mux_o_915;
wire mux_o_916;
wire mux_o_917;
wire mux_o_918;
wire mux_o_919;
wire mux_o_920;
wire mux_o_921;
wire mux_o_922;
wire mux_o_923;
wire mux_o_924;
wire mux_o_925;
wire mux_o_926;
wire mux_o_927;
wire mux_o_928;
wire mux_o_929;
wire mux_o_930;
wire mux_o_931;
wire mux_o_932;
wire mux_o_933;
wire mux_o_934;
wire mux_o_935;
wire mux_o_936;
wire mux_o_937;
wire mux_o_938;
wire mux_o_939;
wire mux_o_940;
wire mux_o_941;
wire mux_o_942;
wire mux_o_943;
wire mux_o_945;
wire mux_o_946;
wire mux_o_947;
wire mux_o_948;
wire mux_o_949;
wire mux_o_950;
wire mux_o_951;
wire mux_o_952;
wire mux_o_953;
wire mux_o_954;
wire mux_o_955;
wire mux_o_956;
wire mux_o_957;
wire mux_o_958;
wire mux_o_959;
wire mux_o_960;
wire mux_o_961;
wire mux_o_962;
wire mux_o_963;
wire mux_o_964;
wire mux_o_965;
wire mux_o_966;
wire mux_o_967;
wire mux_o_968;
wire mux_o_969;
wire mux_o_970;
wire mux_o_971;
wire mux_o_972;
wire mux_o_973;
wire mux_o_974;
wire mux_o_975;
wire mux_o_976;
wire mux_o_977;
wire mux_o_978;
wire mux_o_979;
wire mux_o_980;
wire mux_o_981;
wire mux_o_982;
wire mux_o_983;
wire mux_o_984;
wire mux_o_985;
wire mux_o_986;
wire mux_o_987;
wire mux_o_988;
wire mux_o_989;
wire mux_o_990;
wire mux_o_991;
wire mux_o_992;
wire mux_o_993;
wire mux_o_994;
wire mux_o_995;
wire mux_o_996;
wire mux_o_997;
wire mux_o_998;
wire mux_o_999;
wire mux_o_1000;
wire mux_o_1001;
wire mux_o_1002;
wire mux_o_1003;
wire mux_o_1004;
wire mux_o_1005;
wire mux_o_1006;

ROM16 rom16_inst_0 (
    .DO(rom16_inst_0_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_0.INIT_0 = 16'h0300;

ROM16 rom16_inst_1 (
    .DO(rom16_inst_1_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_1.INIT_0 = 16'h1C27;

ROM16 rom16_inst_2 (
    .DO(rom16_inst_2_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_2.INIT_0 = 16'h1D27;

ROM16 rom16_inst_3 (
    .DO(rom16_inst_3_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_3.INIT_0 = 16'h22B5;

ROM16 rom16_inst_4 (
    .DO(rom16_inst_4_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_4.INIT_0 = 16'h1EB7;

ROM16 rom16_inst_5 (
    .DO(rom16_inst_5_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_5.INIT_0 = 16'h14E3;

ROM16 rom16_inst_6 (
    .DO(rom16_inst_6_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_6.INIT_0 = 16'h3BFC;

ROM16 rom16_inst_7 (
    .DO(rom16_inst_7_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_7.INIT_0 = 16'h2000;

ROM16 rom16_inst_8 (
    .DO(rom16_inst_8_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_8.INIT_0 = 16'h23C9;

ROM16 rom16_inst_9 (
    .DO(rom16_inst_9_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_9.INIT_0 = 16'h2191;

ROM16 rom16_inst_10 (
    .DO(rom16_inst_10_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_10.INIT_0 = 16'h2001;

ROM16 rom16_inst_11 (
    .DO(rom16_inst_11_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_11.INIT_0 = 16'h0001;

ROM16 rom16_inst_12 (
    .DO(rom16_inst_12_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_12.INIT_0 = 16'h0005;

ROM16 rom16_inst_13 (
    .DO(rom16_inst_13_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_13.INIT_0 = 16'h0021;

ROM16 rom16_inst_14 (
    .DO(rom16_inst_14_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_14.INIT_0 = 16'h0003;

ROM16 rom16_inst_15 (
    .DO(rom16_inst_15_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_15.INIT_0 = 16'h1C01;

ROM16 rom16_inst_16 (
    .DO(rom16_inst_16_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_16.INIT_0 = 16'h0000;

ROM16 rom16_inst_17 (
    .DO(rom16_inst_17_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_17.INIT_0 = 16'h0000;

ROM16 rom16_inst_18 (
    .DO(rom16_inst_18_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_18.INIT_0 = 16'h0000;

ROM16 rom16_inst_19 (
    .DO(rom16_inst_19_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_19.INIT_0 = 16'h0000;

ROM16 rom16_inst_20 (
    .DO(rom16_inst_20_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_20.INIT_0 = 16'h0000;

ROM16 rom16_inst_21 (
    .DO(rom16_inst_21_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_21.INIT_0 = 16'h0000;

ROM16 rom16_inst_22 (
    .DO(rom16_inst_22_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_22.INIT_0 = 16'h0000;

ROM16 rom16_inst_23 (
    .DO(rom16_inst_23_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_23.INIT_0 = 16'h0000;

ROM16 rom16_inst_24 (
    .DO(rom16_inst_24_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_24.INIT_0 = 16'h0000;

ROM16 rom16_inst_25 (
    .DO(rom16_inst_25_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_25.INIT_0 = 16'h0000;

ROM16 rom16_inst_26 (
    .DO(rom16_inst_26_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_26.INIT_0 = 16'h0000;

ROM16 rom16_inst_27 (
    .DO(rom16_inst_27_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_27.INIT_0 = 16'h0000;

ROM16 rom16_inst_28 (
    .DO(rom16_inst_28_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_28.INIT_0 = 16'h0000;

ROM16 rom16_inst_29 (
    .DO(rom16_inst_29_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_29.INIT_0 = 16'h0000;

ROM16 rom16_inst_30 (
    .DO(rom16_inst_30_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_30.INIT_0 = 16'h0000;

ROM16 rom16_inst_31 (
    .DO(rom16_inst_31_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_31.INIT_0 = 16'h0000;

ROM16 rom16_inst_32 (
    .DO(rom16_inst_32_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_32.INIT_0 = 16'h0000;

ROM16 rom16_inst_33 (
    .DO(rom16_inst_33_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_33.INIT_0 = 16'h0000;

ROM16 rom16_inst_34 (
    .DO(rom16_inst_34_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_34.INIT_0 = 16'h0000;

ROM16 rom16_inst_35 (
    .DO(rom16_inst_35_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_35.INIT_0 = 16'h0000;

ROM16 rom16_inst_36 (
    .DO(rom16_inst_36_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_36.INIT_0 = 16'h0000;

ROM16 rom16_inst_37 (
    .DO(rom16_inst_37_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_37.INIT_0 = 16'h0000;

ROM16 rom16_inst_38 (
    .DO(rom16_inst_38_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_38.INIT_0 = 16'h0000;

ROM16 rom16_inst_39 (
    .DO(rom16_inst_39_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_39.INIT_0 = 16'h0000;

ROM16 rom16_inst_40 (
    .DO(rom16_inst_40_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_40.INIT_0 = 16'h0000;

ROM16 rom16_inst_41 (
    .DO(rom16_inst_41_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_41.INIT_0 = 16'h0000;

ROM16 rom16_inst_42 (
    .DO(rom16_inst_42_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_42.INIT_0 = 16'h0000;

ROM16 rom16_inst_43 (
    .DO(rom16_inst_43_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_43.INIT_0 = 16'h0000;

ROM16 rom16_inst_44 (
    .DO(rom16_inst_44_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_44.INIT_0 = 16'h0000;

ROM16 rom16_inst_45 (
    .DO(rom16_inst_45_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_45.INIT_0 = 16'h0000;

ROM16 rom16_inst_46 (
    .DO(rom16_inst_46_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_46.INIT_0 = 16'h0000;

ROM16 rom16_inst_47 (
    .DO(rom16_inst_47_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_47.INIT_0 = 16'h0000;

ROM16 rom16_inst_48 (
    .DO(rom16_inst_48_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_48.INIT_0 = 16'h0000;

ROM16 rom16_inst_49 (
    .DO(rom16_inst_49_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_49.INIT_0 = 16'h0000;

ROM16 rom16_inst_50 (
    .DO(rom16_inst_50_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_50.INIT_0 = 16'h0000;

ROM16 rom16_inst_51 (
    .DO(rom16_inst_51_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_51.INIT_0 = 16'h0000;

ROM16 rom16_inst_52 (
    .DO(rom16_inst_52_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_52.INIT_0 = 16'h0000;

ROM16 rom16_inst_53 (
    .DO(rom16_inst_53_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_53.INIT_0 = 16'h0000;

ROM16 rom16_inst_54 (
    .DO(rom16_inst_54_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_54.INIT_0 = 16'h0000;

ROM16 rom16_inst_55 (
    .DO(rom16_inst_55_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_55.INIT_0 = 16'h0000;

ROM16 rom16_inst_56 (
    .DO(rom16_inst_56_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_56.INIT_0 = 16'h0000;

ROM16 rom16_inst_57 (
    .DO(rom16_inst_57_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_57.INIT_0 = 16'h0000;

ROM16 rom16_inst_58 (
    .DO(rom16_inst_58_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_58.INIT_0 = 16'h0000;

ROM16 rom16_inst_59 (
    .DO(rom16_inst_59_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_59.INIT_0 = 16'h0000;

ROM16 rom16_inst_60 (
    .DO(rom16_inst_60_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_60.INIT_0 = 16'h0000;

ROM16 rom16_inst_61 (
    .DO(rom16_inst_61_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_61.INIT_0 = 16'h0000;

ROM16 rom16_inst_62 (
    .DO(rom16_inst_62_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_62.INIT_0 = 16'h0000;

ROM16 rom16_inst_63 (
    .DO(rom16_inst_63_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_63.INIT_0 = 16'h0000;

ROM16 rom16_inst_64 (
    .DO(rom16_inst_64_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_64.INIT_0 = 16'h0000;

ROM16 rom16_inst_65 (
    .DO(rom16_inst_65_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_65.INIT_0 = 16'h0000;

ROM16 rom16_inst_66 (
    .DO(rom16_inst_66_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_66.INIT_0 = 16'h0000;

ROM16 rom16_inst_67 (
    .DO(rom16_inst_67_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_67.INIT_0 = 16'h0000;

ROM16 rom16_inst_68 (
    .DO(rom16_inst_68_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_68.INIT_0 = 16'h0000;

ROM16 rom16_inst_69 (
    .DO(rom16_inst_69_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_69.INIT_0 = 16'h0000;

ROM16 rom16_inst_70 (
    .DO(rom16_inst_70_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_70.INIT_0 = 16'h0000;

ROM16 rom16_inst_71 (
    .DO(rom16_inst_71_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_71.INIT_0 = 16'h0000;

ROM16 rom16_inst_72 (
    .DO(rom16_inst_72_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_72.INIT_0 = 16'h0000;

ROM16 rom16_inst_73 (
    .DO(rom16_inst_73_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_73.INIT_0 = 16'h0000;

ROM16 rom16_inst_74 (
    .DO(rom16_inst_74_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_74.INIT_0 = 16'h0000;

ROM16 rom16_inst_75 (
    .DO(rom16_inst_75_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_75.INIT_0 = 16'h0000;

ROM16 rom16_inst_76 (
    .DO(rom16_inst_76_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_76.INIT_0 = 16'h0000;

ROM16 rom16_inst_77 (
    .DO(rom16_inst_77_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_77.INIT_0 = 16'h0000;

ROM16 rom16_inst_78 (
    .DO(rom16_inst_78_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_78.INIT_0 = 16'h0000;

ROM16 rom16_inst_79 (
    .DO(rom16_inst_79_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_79.INIT_0 = 16'h0000;

ROM16 rom16_inst_80 (
    .DO(rom16_inst_80_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_80.INIT_0 = 16'h0000;

ROM16 rom16_inst_81 (
    .DO(rom16_inst_81_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_81.INIT_0 = 16'h0000;

ROM16 rom16_inst_82 (
    .DO(rom16_inst_82_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_82.INIT_0 = 16'h0000;

ROM16 rom16_inst_83 (
    .DO(rom16_inst_83_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_83.INIT_0 = 16'h0000;

ROM16 rom16_inst_84 (
    .DO(rom16_inst_84_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_84.INIT_0 = 16'h0000;

ROM16 rom16_inst_85 (
    .DO(rom16_inst_85_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_85.INIT_0 = 16'h0000;

ROM16 rom16_inst_86 (
    .DO(rom16_inst_86_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_86.INIT_0 = 16'h0000;

ROM16 rom16_inst_87 (
    .DO(rom16_inst_87_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_87.INIT_0 = 16'h0000;

ROM16 rom16_inst_88 (
    .DO(rom16_inst_88_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_88.INIT_0 = 16'h0000;

ROM16 rom16_inst_89 (
    .DO(rom16_inst_89_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_89.INIT_0 = 16'h0000;

ROM16 rom16_inst_90 (
    .DO(rom16_inst_90_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_90.INIT_0 = 16'h0000;

ROM16 rom16_inst_91 (
    .DO(rom16_inst_91_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_91.INIT_0 = 16'h0000;

ROM16 rom16_inst_92 (
    .DO(rom16_inst_92_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_92.INIT_0 = 16'h0000;

ROM16 rom16_inst_93 (
    .DO(rom16_inst_93_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_93.INIT_0 = 16'h0000;

ROM16 rom16_inst_94 (
    .DO(rom16_inst_94_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_94.INIT_0 = 16'h0000;

ROM16 rom16_inst_95 (
    .DO(rom16_inst_95_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_95.INIT_0 = 16'h0000;

ROM16 rom16_inst_96 (
    .DO(rom16_inst_96_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_96.INIT_0 = 16'h0000;

ROM16 rom16_inst_97 (
    .DO(rom16_inst_97_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_97.INIT_0 = 16'h0000;

ROM16 rom16_inst_98 (
    .DO(rom16_inst_98_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_98.INIT_0 = 16'h0000;

ROM16 rom16_inst_99 (
    .DO(rom16_inst_99_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_99.INIT_0 = 16'h0000;

ROM16 rom16_inst_100 (
    .DO(rom16_inst_100_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_100.INIT_0 = 16'h0000;

ROM16 rom16_inst_101 (
    .DO(rom16_inst_101_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_101.INIT_0 = 16'h0000;

ROM16 rom16_inst_102 (
    .DO(rom16_inst_102_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_102.INIT_0 = 16'h0000;

ROM16 rom16_inst_103 (
    .DO(rom16_inst_103_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_103.INIT_0 = 16'h0000;

ROM16 rom16_inst_104 (
    .DO(rom16_inst_104_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_104.INIT_0 = 16'h0000;

ROM16 rom16_inst_105 (
    .DO(rom16_inst_105_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_105.INIT_0 = 16'h0000;

ROM16 rom16_inst_106 (
    .DO(rom16_inst_106_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_106.INIT_0 = 16'h0000;

ROM16 rom16_inst_107 (
    .DO(rom16_inst_107_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_107.INIT_0 = 16'h0000;

ROM16 rom16_inst_108 (
    .DO(rom16_inst_108_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_108.INIT_0 = 16'h0000;

ROM16 rom16_inst_109 (
    .DO(rom16_inst_109_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_109.INIT_0 = 16'h0000;

ROM16 rom16_inst_110 (
    .DO(rom16_inst_110_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_110.INIT_0 = 16'h0000;

ROM16 rom16_inst_111 (
    .DO(rom16_inst_111_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_111.INIT_0 = 16'h0000;

ROM16 rom16_inst_112 (
    .DO(rom16_inst_112_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_112.INIT_0 = 16'h0000;

ROM16 rom16_inst_113 (
    .DO(rom16_inst_113_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_113.INIT_0 = 16'h0000;

ROM16 rom16_inst_114 (
    .DO(rom16_inst_114_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_114.INIT_0 = 16'h0000;

ROM16 rom16_inst_115 (
    .DO(rom16_inst_115_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_115.INIT_0 = 16'h0000;

ROM16 rom16_inst_116 (
    .DO(rom16_inst_116_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_116.INIT_0 = 16'h0000;

ROM16 rom16_inst_117 (
    .DO(rom16_inst_117_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_117.INIT_0 = 16'h0000;

ROM16 rom16_inst_118 (
    .DO(rom16_inst_118_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_118.INIT_0 = 16'h0000;

ROM16 rom16_inst_119 (
    .DO(rom16_inst_119_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_119.INIT_0 = 16'h0000;

ROM16 rom16_inst_120 (
    .DO(rom16_inst_120_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_120.INIT_0 = 16'h0000;

ROM16 rom16_inst_121 (
    .DO(rom16_inst_121_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_121.INIT_0 = 16'h0000;

ROM16 rom16_inst_122 (
    .DO(rom16_inst_122_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_122.INIT_0 = 16'h0000;

ROM16 rom16_inst_123 (
    .DO(rom16_inst_123_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_123.INIT_0 = 16'h0000;

ROM16 rom16_inst_124 (
    .DO(rom16_inst_124_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_124.INIT_0 = 16'h0000;

ROM16 rom16_inst_125 (
    .DO(rom16_inst_125_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_125.INIT_0 = 16'h0000;

ROM16 rom16_inst_126 (
    .DO(rom16_inst_126_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_126.INIT_0 = 16'h0000;

ROM16 rom16_inst_127 (
    .DO(rom16_inst_127_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_127.INIT_0 = 16'h0000;

ROM16 rom16_inst_128 (
    .DO(rom16_inst_128_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_128.INIT_0 = 16'h0000;

ROM16 rom16_inst_129 (
    .DO(rom16_inst_129_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_129.INIT_0 = 16'h0000;

ROM16 rom16_inst_130 (
    .DO(rom16_inst_130_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_130.INIT_0 = 16'h0000;

ROM16 rom16_inst_131 (
    .DO(rom16_inst_131_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_131.INIT_0 = 16'h0000;

ROM16 rom16_inst_132 (
    .DO(rom16_inst_132_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_132.INIT_0 = 16'h0000;

ROM16 rom16_inst_133 (
    .DO(rom16_inst_133_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_133.INIT_0 = 16'h0000;

ROM16 rom16_inst_134 (
    .DO(rom16_inst_134_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_134.INIT_0 = 16'h0000;

ROM16 rom16_inst_135 (
    .DO(rom16_inst_135_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_135.INIT_0 = 16'h0000;

ROM16 rom16_inst_136 (
    .DO(rom16_inst_136_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_136.INIT_0 = 16'h0000;

ROM16 rom16_inst_137 (
    .DO(rom16_inst_137_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_137.INIT_0 = 16'h0000;

ROM16 rom16_inst_138 (
    .DO(rom16_inst_138_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_138.INIT_0 = 16'h0000;

ROM16 rom16_inst_139 (
    .DO(rom16_inst_139_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_139.INIT_0 = 16'h0000;

ROM16 rom16_inst_140 (
    .DO(rom16_inst_140_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_140.INIT_0 = 16'h0000;

ROM16 rom16_inst_141 (
    .DO(rom16_inst_141_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_141.INIT_0 = 16'h0000;

ROM16 rom16_inst_142 (
    .DO(rom16_inst_142_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_142.INIT_0 = 16'h0000;

ROM16 rom16_inst_143 (
    .DO(rom16_inst_143_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_143.INIT_0 = 16'h0000;

ROM16 rom16_inst_144 (
    .DO(rom16_inst_144_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_144.INIT_0 = 16'h0000;

ROM16 rom16_inst_145 (
    .DO(rom16_inst_145_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_145.INIT_0 = 16'h0000;

ROM16 rom16_inst_146 (
    .DO(rom16_inst_146_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_146.INIT_0 = 16'h0000;

ROM16 rom16_inst_147 (
    .DO(rom16_inst_147_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_147.INIT_0 = 16'h0000;

ROM16 rom16_inst_148 (
    .DO(rom16_inst_148_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_148.INIT_0 = 16'h0000;

ROM16 rom16_inst_149 (
    .DO(rom16_inst_149_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_149.INIT_0 = 16'h0000;

ROM16 rom16_inst_150 (
    .DO(rom16_inst_150_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_150.INIT_0 = 16'h0000;

ROM16 rom16_inst_151 (
    .DO(rom16_inst_151_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_151.INIT_0 = 16'h0000;

ROM16 rom16_inst_152 (
    .DO(rom16_inst_152_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_152.INIT_0 = 16'h0000;

ROM16 rom16_inst_153 (
    .DO(rom16_inst_153_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_153.INIT_0 = 16'h0000;

ROM16 rom16_inst_154 (
    .DO(rom16_inst_154_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_154.INIT_0 = 16'h0000;

ROM16 rom16_inst_155 (
    .DO(rom16_inst_155_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_155.INIT_0 = 16'h0000;

ROM16 rom16_inst_156 (
    .DO(rom16_inst_156_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_156.INIT_0 = 16'h0000;

ROM16 rom16_inst_157 (
    .DO(rom16_inst_157_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_157.INIT_0 = 16'h0000;

ROM16 rom16_inst_158 (
    .DO(rom16_inst_158_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_158.INIT_0 = 16'h0000;

ROM16 rom16_inst_159 (
    .DO(rom16_inst_159_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_159.INIT_0 = 16'h0000;

ROM16 rom16_inst_160 (
    .DO(rom16_inst_160_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_160.INIT_0 = 16'h0000;

ROM16 rom16_inst_161 (
    .DO(rom16_inst_161_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_161.INIT_0 = 16'h0000;

ROM16 rom16_inst_162 (
    .DO(rom16_inst_162_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_162.INIT_0 = 16'h0000;

ROM16 rom16_inst_163 (
    .DO(rom16_inst_163_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_163.INIT_0 = 16'h0000;

ROM16 rom16_inst_164 (
    .DO(rom16_inst_164_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_164.INIT_0 = 16'h0000;

ROM16 rom16_inst_165 (
    .DO(rom16_inst_165_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_165.INIT_0 = 16'h0000;

ROM16 rom16_inst_166 (
    .DO(rom16_inst_166_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_166.INIT_0 = 16'h0000;

ROM16 rom16_inst_167 (
    .DO(rom16_inst_167_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_167.INIT_0 = 16'h0000;

ROM16 rom16_inst_168 (
    .DO(rom16_inst_168_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_168.INIT_0 = 16'h0000;

ROM16 rom16_inst_169 (
    .DO(rom16_inst_169_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_169.INIT_0 = 16'h0000;

ROM16 rom16_inst_170 (
    .DO(rom16_inst_170_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_170.INIT_0 = 16'h0000;

ROM16 rom16_inst_171 (
    .DO(rom16_inst_171_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_171.INIT_0 = 16'h0000;

ROM16 rom16_inst_172 (
    .DO(rom16_inst_172_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_172.INIT_0 = 16'h0000;

ROM16 rom16_inst_173 (
    .DO(rom16_inst_173_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_173.INIT_0 = 16'h0000;

ROM16 rom16_inst_174 (
    .DO(rom16_inst_174_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_174.INIT_0 = 16'h0000;

ROM16 rom16_inst_175 (
    .DO(rom16_inst_175_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_175.INIT_0 = 16'h0000;

ROM16 rom16_inst_176 (
    .DO(rom16_inst_176_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_176.INIT_0 = 16'h0000;

ROM16 rom16_inst_177 (
    .DO(rom16_inst_177_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_177.INIT_0 = 16'h0000;

ROM16 rom16_inst_178 (
    .DO(rom16_inst_178_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_178.INIT_0 = 16'h0000;

ROM16 rom16_inst_179 (
    .DO(rom16_inst_179_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_179.INIT_0 = 16'h0000;

ROM16 rom16_inst_180 (
    .DO(rom16_inst_180_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_180.INIT_0 = 16'h0000;

ROM16 rom16_inst_181 (
    .DO(rom16_inst_181_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_181.INIT_0 = 16'h0000;

ROM16 rom16_inst_182 (
    .DO(rom16_inst_182_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_182.INIT_0 = 16'h0000;

ROM16 rom16_inst_183 (
    .DO(rom16_inst_183_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_183.INIT_0 = 16'h0000;

ROM16 rom16_inst_184 (
    .DO(rom16_inst_184_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_184.INIT_0 = 16'h0000;

ROM16 rom16_inst_185 (
    .DO(rom16_inst_185_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_185.INIT_0 = 16'h0000;

ROM16 rom16_inst_186 (
    .DO(rom16_inst_186_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_186.INIT_0 = 16'h0000;

ROM16 rom16_inst_187 (
    .DO(rom16_inst_187_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_187.INIT_0 = 16'h0000;

ROM16 rom16_inst_188 (
    .DO(rom16_inst_188_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_188.INIT_0 = 16'h0000;

ROM16 rom16_inst_189 (
    .DO(rom16_inst_189_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_189.INIT_0 = 16'h0000;

ROM16 rom16_inst_190 (
    .DO(rom16_inst_190_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_190.INIT_0 = 16'h0000;

ROM16 rom16_inst_191 (
    .DO(rom16_inst_191_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_191.INIT_0 = 16'h0000;

ROM16 rom16_inst_192 (
    .DO(rom16_inst_192_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_192.INIT_0 = 16'h0000;

ROM16 rom16_inst_193 (
    .DO(rom16_inst_193_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_193.INIT_0 = 16'h0000;

ROM16 rom16_inst_194 (
    .DO(rom16_inst_194_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_194.INIT_0 = 16'h0000;

ROM16 rom16_inst_195 (
    .DO(rom16_inst_195_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_195.INIT_0 = 16'h0000;

ROM16 rom16_inst_196 (
    .DO(rom16_inst_196_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_196.INIT_0 = 16'h0000;

ROM16 rom16_inst_197 (
    .DO(rom16_inst_197_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_197.INIT_0 = 16'h0000;

ROM16 rom16_inst_198 (
    .DO(rom16_inst_198_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_198.INIT_0 = 16'h0000;

ROM16 rom16_inst_199 (
    .DO(rom16_inst_199_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_199.INIT_0 = 16'h0000;

ROM16 rom16_inst_200 (
    .DO(rom16_inst_200_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_200.INIT_0 = 16'h0000;

ROM16 rom16_inst_201 (
    .DO(rom16_inst_201_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_201.INIT_0 = 16'h0000;

ROM16 rom16_inst_202 (
    .DO(rom16_inst_202_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_202.INIT_0 = 16'h0000;

ROM16 rom16_inst_203 (
    .DO(rom16_inst_203_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_203.INIT_0 = 16'h0000;

ROM16 rom16_inst_204 (
    .DO(rom16_inst_204_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_204.INIT_0 = 16'h0000;

ROM16 rom16_inst_205 (
    .DO(rom16_inst_205_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_205.INIT_0 = 16'h0000;

ROM16 rom16_inst_206 (
    .DO(rom16_inst_206_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_206.INIT_0 = 16'h0000;

ROM16 rom16_inst_207 (
    .DO(rom16_inst_207_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_207.INIT_0 = 16'h0000;

ROM16 rom16_inst_208 (
    .DO(rom16_inst_208_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_208.INIT_0 = 16'h0000;

ROM16 rom16_inst_209 (
    .DO(rom16_inst_209_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_209.INIT_0 = 16'h0000;

ROM16 rom16_inst_210 (
    .DO(rom16_inst_210_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_210.INIT_0 = 16'h0000;

ROM16 rom16_inst_211 (
    .DO(rom16_inst_211_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_211.INIT_0 = 16'h0000;

ROM16 rom16_inst_212 (
    .DO(rom16_inst_212_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_212.INIT_0 = 16'h0000;

ROM16 rom16_inst_213 (
    .DO(rom16_inst_213_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_213.INIT_0 = 16'h0000;

ROM16 rom16_inst_214 (
    .DO(rom16_inst_214_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_214.INIT_0 = 16'h0000;

ROM16 rom16_inst_215 (
    .DO(rom16_inst_215_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_215.INIT_0 = 16'h0000;

ROM16 rom16_inst_216 (
    .DO(rom16_inst_216_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_216.INIT_0 = 16'h0000;

ROM16 rom16_inst_217 (
    .DO(rom16_inst_217_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_217.INIT_0 = 16'h0000;

ROM16 rom16_inst_218 (
    .DO(rom16_inst_218_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_218.INIT_0 = 16'h0000;

ROM16 rom16_inst_219 (
    .DO(rom16_inst_219_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_219.INIT_0 = 16'h0000;

ROM16 rom16_inst_220 (
    .DO(rom16_inst_220_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_220.INIT_0 = 16'h0000;

ROM16 rom16_inst_221 (
    .DO(rom16_inst_221_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_221.INIT_0 = 16'h0000;

ROM16 rom16_inst_222 (
    .DO(rom16_inst_222_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_222.INIT_0 = 16'h0000;

ROM16 rom16_inst_223 (
    .DO(rom16_inst_223_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_223.INIT_0 = 16'h0000;

ROM16 rom16_inst_224 (
    .DO(rom16_inst_224_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_224.INIT_0 = 16'h0000;

ROM16 rom16_inst_225 (
    .DO(rom16_inst_225_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_225.INIT_0 = 16'h0000;

ROM16 rom16_inst_226 (
    .DO(rom16_inst_226_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_226.INIT_0 = 16'h0000;

ROM16 rom16_inst_227 (
    .DO(rom16_inst_227_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_227.INIT_0 = 16'h0000;

ROM16 rom16_inst_228 (
    .DO(rom16_inst_228_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_228.INIT_0 = 16'h0000;

ROM16 rom16_inst_229 (
    .DO(rom16_inst_229_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_229.INIT_0 = 16'h0000;

ROM16 rom16_inst_230 (
    .DO(rom16_inst_230_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_230.INIT_0 = 16'h0000;

ROM16 rom16_inst_231 (
    .DO(rom16_inst_231_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_231.INIT_0 = 16'h0000;

ROM16 rom16_inst_232 (
    .DO(rom16_inst_232_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_232.INIT_0 = 16'h0000;

ROM16 rom16_inst_233 (
    .DO(rom16_inst_233_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_233.INIT_0 = 16'h0000;

ROM16 rom16_inst_234 (
    .DO(rom16_inst_234_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_234.INIT_0 = 16'h0000;

ROM16 rom16_inst_235 (
    .DO(rom16_inst_235_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_235.INIT_0 = 16'h0000;

ROM16 rom16_inst_236 (
    .DO(rom16_inst_236_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_236.INIT_0 = 16'h0000;

ROM16 rom16_inst_237 (
    .DO(rom16_inst_237_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_237.INIT_0 = 16'h0000;

ROM16 rom16_inst_238 (
    .DO(rom16_inst_238_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_238.INIT_0 = 16'h0000;

ROM16 rom16_inst_239 (
    .DO(rom16_inst_239_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_239.INIT_0 = 16'h0000;

ROM16 rom16_inst_240 (
    .DO(rom16_inst_240_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_240.INIT_0 = 16'h0000;

ROM16 rom16_inst_241 (
    .DO(rom16_inst_241_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_241.INIT_0 = 16'h0000;

ROM16 rom16_inst_242 (
    .DO(rom16_inst_242_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_242.INIT_0 = 16'h0000;

ROM16 rom16_inst_243 (
    .DO(rom16_inst_243_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_243.INIT_0 = 16'h0000;

ROM16 rom16_inst_244 (
    .DO(rom16_inst_244_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_244.INIT_0 = 16'h0000;

ROM16 rom16_inst_245 (
    .DO(rom16_inst_245_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_245.INIT_0 = 16'h0000;

ROM16 rom16_inst_246 (
    .DO(rom16_inst_246_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_246.INIT_0 = 16'h0000;

ROM16 rom16_inst_247 (
    .DO(rom16_inst_247_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_247.INIT_0 = 16'h0000;

ROM16 rom16_inst_248 (
    .DO(rom16_inst_248_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_248.INIT_0 = 16'h0000;

ROM16 rom16_inst_249 (
    .DO(rom16_inst_249_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_249.INIT_0 = 16'h0000;

ROM16 rom16_inst_250 (
    .DO(rom16_inst_250_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_250.INIT_0 = 16'h0000;

ROM16 rom16_inst_251 (
    .DO(rom16_inst_251_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_251.INIT_0 = 16'h0000;

ROM16 rom16_inst_252 (
    .DO(rom16_inst_252_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_252.INIT_0 = 16'h0000;

ROM16 rom16_inst_253 (
    .DO(rom16_inst_253_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_253.INIT_0 = 16'h0000;

ROM16 rom16_inst_254 (
    .DO(rom16_inst_254_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_254.INIT_0 = 16'h0000;

ROM16 rom16_inst_255 (
    .DO(rom16_inst_255_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_255.INIT_0 = 16'h0000;

ROM16 rom16_inst_256 (
    .DO(rom16_inst_256_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_256.INIT_0 = 16'h0000;

ROM16 rom16_inst_257 (
    .DO(rom16_inst_257_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_257.INIT_0 = 16'h0000;

ROM16 rom16_inst_258 (
    .DO(rom16_inst_258_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_258.INIT_0 = 16'h0000;

ROM16 rom16_inst_259 (
    .DO(rom16_inst_259_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_259.INIT_0 = 16'h0000;

ROM16 rom16_inst_260 (
    .DO(rom16_inst_260_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_260.INIT_0 = 16'h0000;

ROM16 rom16_inst_261 (
    .DO(rom16_inst_261_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_261.INIT_0 = 16'h0000;

ROM16 rom16_inst_262 (
    .DO(rom16_inst_262_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_262.INIT_0 = 16'h0000;

ROM16 rom16_inst_263 (
    .DO(rom16_inst_263_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_263.INIT_0 = 16'h0000;

ROM16 rom16_inst_264 (
    .DO(rom16_inst_264_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_264.INIT_0 = 16'h0000;

ROM16 rom16_inst_265 (
    .DO(rom16_inst_265_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_265.INIT_0 = 16'h0000;

ROM16 rom16_inst_266 (
    .DO(rom16_inst_266_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_266.INIT_0 = 16'h0000;

ROM16 rom16_inst_267 (
    .DO(rom16_inst_267_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_267.INIT_0 = 16'h0000;

ROM16 rom16_inst_268 (
    .DO(rom16_inst_268_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_268.INIT_0 = 16'h0000;

ROM16 rom16_inst_269 (
    .DO(rom16_inst_269_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_269.INIT_0 = 16'h0000;

ROM16 rom16_inst_270 (
    .DO(rom16_inst_270_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_270.INIT_0 = 16'h0000;

ROM16 rom16_inst_271 (
    .DO(rom16_inst_271_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_271.INIT_0 = 16'h0000;

ROM16 rom16_inst_272 (
    .DO(rom16_inst_272_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_272.INIT_0 = 16'h0000;

ROM16 rom16_inst_273 (
    .DO(rom16_inst_273_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_273.INIT_0 = 16'h0000;

ROM16 rom16_inst_274 (
    .DO(rom16_inst_274_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_274.INIT_0 = 16'h0000;

ROM16 rom16_inst_275 (
    .DO(rom16_inst_275_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_275.INIT_0 = 16'h0000;

ROM16 rom16_inst_276 (
    .DO(rom16_inst_276_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_276.INIT_0 = 16'h0000;

ROM16 rom16_inst_277 (
    .DO(rom16_inst_277_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_277.INIT_0 = 16'h0000;

ROM16 rom16_inst_278 (
    .DO(rom16_inst_278_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_278.INIT_0 = 16'h0000;

ROM16 rom16_inst_279 (
    .DO(rom16_inst_279_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_279.INIT_0 = 16'h0000;

ROM16 rom16_inst_280 (
    .DO(rom16_inst_280_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_280.INIT_0 = 16'h0000;

ROM16 rom16_inst_281 (
    .DO(rom16_inst_281_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_281.INIT_0 = 16'h0000;

ROM16 rom16_inst_282 (
    .DO(rom16_inst_282_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_282.INIT_0 = 16'h0000;

ROM16 rom16_inst_283 (
    .DO(rom16_inst_283_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_283.INIT_0 = 16'h0000;

ROM16 rom16_inst_284 (
    .DO(rom16_inst_284_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_284.INIT_0 = 16'h0000;

ROM16 rom16_inst_285 (
    .DO(rom16_inst_285_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_285.INIT_0 = 16'h0000;

ROM16 rom16_inst_286 (
    .DO(rom16_inst_286_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_286.INIT_0 = 16'h0000;

ROM16 rom16_inst_287 (
    .DO(rom16_inst_287_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_287.INIT_0 = 16'h0000;

ROM16 rom16_inst_288 (
    .DO(rom16_inst_288_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_288.INIT_0 = 16'h0000;

ROM16 rom16_inst_289 (
    .DO(rom16_inst_289_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_289.INIT_0 = 16'h0000;

ROM16 rom16_inst_290 (
    .DO(rom16_inst_290_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_290.INIT_0 = 16'h0000;

ROM16 rom16_inst_291 (
    .DO(rom16_inst_291_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_291.INIT_0 = 16'h0000;

ROM16 rom16_inst_292 (
    .DO(rom16_inst_292_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_292.INIT_0 = 16'h0000;

ROM16 rom16_inst_293 (
    .DO(rom16_inst_293_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_293.INIT_0 = 16'h0000;

ROM16 rom16_inst_294 (
    .DO(rom16_inst_294_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_294.INIT_0 = 16'h0000;

ROM16 rom16_inst_295 (
    .DO(rom16_inst_295_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_295.INIT_0 = 16'h0000;

ROM16 rom16_inst_296 (
    .DO(rom16_inst_296_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_296.INIT_0 = 16'h0000;

ROM16 rom16_inst_297 (
    .DO(rom16_inst_297_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_297.INIT_0 = 16'h0000;

ROM16 rom16_inst_298 (
    .DO(rom16_inst_298_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_298.INIT_0 = 16'h0000;

ROM16 rom16_inst_299 (
    .DO(rom16_inst_299_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_299.INIT_0 = 16'h0000;

ROM16 rom16_inst_300 (
    .DO(rom16_inst_300_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_300.INIT_0 = 16'h0000;

ROM16 rom16_inst_301 (
    .DO(rom16_inst_301_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_301.INIT_0 = 16'h0000;

ROM16 rom16_inst_302 (
    .DO(rom16_inst_302_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_302.INIT_0 = 16'h0000;

ROM16 rom16_inst_303 (
    .DO(rom16_inst_303_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_303.INIT_0 = 16'h0000;

ROM16 rom16_inst_304 (
    .DO(rom16_inst_304_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_304.INIT_0 = 16'h0000;

ROM16 rom16_inst_305 (
    .DO(rom16_inst_305_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_305.INIT_0 = 16'h0000;

ROM16 rom16_inst_306 (
    .DO(rom16_inst_306_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_306.INIT_0 = 16'h0000;

ROM16 rom16_inst_307 (
    .DO(rom16_inst_307_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_307.INIT_0 = 16'h0000;

ROM16 rom16_inst_308 (
    .DO(rom16_inst_308_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_308.INIT_0 = 16'h0000;

ROM16 rom16_inst_309 (
    .DO(rom16_inst_309_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_309.INIT_0 = 16'h0000;

ROM16 rom16_inst_310 (
    .DO(rom16_inst_310_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_310.INIT_0 = 16'h0000;

ROM16 rom16_inst_311 (
    .DO(rom16_inst_311_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_311.INIT_0 = 16'h0000;

ROM16 rom16_inst_312 (
    .DO(rom16_inst_312_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_312.INIT_0 = 16'h0000;

ROM16 rom16_inst_313 (
    .DO(rom16_inst_313_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_313.INIT_0 = 16'h0000;

ROM16 rom16_inst_314 (
    .DO(rom16_inst_314_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_314.INIT_0 = 16'h0000;

ROM16 rom16_inst_315 (
    .DO(rom16_inst_315_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_315.INIT_0 = 16'h0000;

ROM16 rom16_inst_316 (
    .DO(rom16_inst_316_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_316.INIT_0 = 16'h0000;

ROM16 rom16_inst_317 (
    .DO(rom16_inst_317_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_317.INIT_0 = 16'h0000;

ROM16 rom16_inst_318 (
    .DO(rom16_inst_318_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_318.INIT_0 = 16'h0000;

ROM16 rom16_inst_319 (
    .DO(rom16_inst_319_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_319.INIT_0 = 16'h0000;

ROM16 rom16_inst_320 (
    .DO(rom16_inst_320_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_320.INIT_0 = 16'h0000;

ROM16 rom16_inst_321 (
    .DO(rom16_inst_321_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_321.INIT_0 = 16'h0000;

ROM16 rom16_inst_322 (
    .DO(rom16_inst_322_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_322.INIT_0 = 16'h0000;

ROM16 rom16_inst_323 (
    .DO(rom16_inst_323_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_323.INIT_0 = 16'h0000;

ROM16 rom16_inst_324 (
    .DO(rom16_inst_324_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_324.INIT_0 = 16'h0000;

ROM16 rom16_inst_325 (
    .DO(rom16_inst_325_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_325.INIT_0 = 16'h0000;

ROM16 rom16_inst_326 (
    .DO(rom16_inst_326_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_326.INIT_0 = 16'h0000;

ROM16 rom16_inst_327 (
    .DO(rom16_inst_327_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_327.INIT_0 = 16'h0000;

ROM16 rom16_inst_328 (
    .DO(rom16_inst_328_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_328.INIT_0 = 16'h0000;

ROM16 rom16_inst_329 (
    .DO(rom16_inst_329_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_329.INIT_0 = 16'h0000;

ROM16 rom16_inst_330 (
    .DO(rom16_inst_330_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_330.INIT_0 = 16'h0000;

ROM16 rom16_inst_331 (
    .DO(rom16_inst_331_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_331.INIT_0 = 16'h0000;

ROM16 rom16_inst_332 (
    .DO(rom16_inst_332_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_332.INIT_0 = 16'h0000;

ROM16 rom16_inst_333 (
    .DO(rom16_inst_333_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_333.INIT_0 = 16'h0000;

ROM16 rom16_inst_334 (
    .DO(rom16_inst_334_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_334.INIT_0 = 16'h0000;

ROM16 rom16_inst_335 (
    .DO(rom16_inst_335_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_335.INIT_0 = 16'h0000;

ROM16 rom16_inst_336 (
    .DO(rom16_inst_336_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_336.INIT_0 = 16'h0000;

ROM16 rom16_inst_337 (
    .DO(rom16_inst_337_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_337.INIT_0 = 16'h0000;

ROM16 rom16_inst_338 (
    .DO(rom16_inst_338_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_338.INIT_0 = 16'h0000;

ROM16 rom16_inst_339 (
    .DO(rom16_inst_339_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_339.INIT_0 = 16'h0000;

ROM16 rom16_inst_340 (
    .DO(rom16_inst_340_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_340.INIT_0 = 16'h0000;

ROM16 rom16_inst_341 (
    .DO(rom16_inst_341_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_341.INIT_0 = 16'h0000;

ROM16 rom16_inst_342 (
    .DO(rom16_inst_342_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_342.INIT_0 = 16'h0000;

ROM16 rom16_inst_343 (
    .DO(rom16_inst_343_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_343.INIT_0 = 16'h0000;

ROM16 rom16_inst_344 (
    .DO(rom16_inst_344_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_344.INIT_0 = 16'h0000;

ROM16 rom16_inst_345 (
    .DO(rom16_inst_345_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_345.INIT_0 = 16'h0000;

ROM16 rom16_inst_346 (
    .DO(rom16_inst_346_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_346.INIT_0 = 16'h0000;

ROM16 rom16_inst_347 (
    .DO(rom16_inst_347_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_347.INIT_0 = 16'h0000;

ROM16 rom16_inst_348 (
    .DO(rom16_inst_348_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_348.INIT_0 = 16'h0000;

ROM16 rom16_inst_349 (
    .DO(rom16_inst_349_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_349.INIT_0 = 16'h0000;

ROM16 rom16_inst_350 (
    .DO(rom16_inst_350_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_350.INIT_0 = 16'h0000;

ROM16 rom16_inst_351 (
    .DO(rom16_inst_351_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_351.INIT_0 = 16'h0000;

ROM16 rom16_inst_352 (
    .DO(rom16_inst_352_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_352.INIT_0 = 16'h0000;

ROM16 rom16_inst_353 (
    .DO(rom16_inst_353_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_353.INIT_0 = 16'h0000;

ROM16 rom16_inst_354 (
    .DO(rom16_inst_354_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_354.INIT_0 = 16'h0000;

ROM16 rom16_inst_355 (
    .DO(rom16_inst_355_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_355.INIT_0 = 16'h0000;

ROM16 rom16_inst_356 (
    .DO(rom16_inst_356_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_356.INIT_0 = 16'h0000;

ROM16 rom16_inst_357 (
    .DO(rom16_inst_357_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_357.INIT_0 = 16'h0000;

ROM16 rom16_inst_358 (
    .DO(rom16_inst_358_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_358.INIT_0 = 16'h0000;

ROM16 rom16_inst_359 (
    .DO(rom16_inst_359_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_359.INIT_0 = 16'h0000;

ROM16 rom16_inst_360 (
    .DO(rom16_inst_360_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_360.INIT_0 = 16'h0000;

ROM16 rom16_inst_361 (
    .DO(rom16_inst_361_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_361.INIT_0 = 16'h0000;

ROM16 rom16_inst_362 (
    .DO(rom16_inst_362_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_362.INIT_0 = 16'h0000;

ROM16 rom16_inst_363 (
    .DO(rom16_inst_363_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_363.INIT_0 = 16'h0000;

ROM16 rom16_inst_364 (
    .DO(rom16_inst_364_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_364.INIT_0 = 16'h0000;

ROM16 rom16_inst_365 (
    .DO(rom16_inst_365_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_365.INIT_0 = 16'h0000;

ROM16 rom16_inst_366 (
    .DO(rom16_inst_366_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_366.INIT_0 = 16'h0000;

ROM16 rom16_inst_367 (
    .DO(rom16_inst_367_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_367.INIT_0 = 16'h0000;

ROM16 rom16_inst_368 (
    .DO(rom16_inst_368_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_368.INIT_0 = 16'h0000;

ROM16 rom16_inst_369 (
    .DO(rom16_inst_369_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_369.INIT_0 = 16'h0000;

ROM16 rom16_inst_370 (
    .DO(rom16_inst_370_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_370.INIT_0 = 16'h0000;

ROM16 rom16_inst_371 (
    .DO(rom16_inst_371_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_371.INIT_0 = 16'h0000;

ROM16 rom16_inst_372 (
    .DO(rom16_inst_372_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_372.INIT_0 = 16'h0000;

ROM16 rom16_inst_373 (
    .DO(rom16_inst_373_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_373.INIT_0 = 16'h0000;

ROM16 rom16_inst_374 (
    .DO(rom16_inst_374_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_374.INIT_0 = 16'h0000;

ROM16 rom16_inst_375 (
    .DO(rom16_inst_375_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_375.INIT_0 = 16'h0000;

ROM16 rom16_inst_376 (
    .DO(rom16_inst_376_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_376.INIT_0 = 16'h0000;

ROM16 rom16_inst_377 (
    .DO(rom16_inst_377_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_377.INIT_0 = 16'h0000;

ROM16 rom16_inst_378 (
    .DO(rom16_inst_378_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_378.INIT_0 = 16'h0000;

ROM16 rom16_inst_379 (
    .DO(rom16_inst_379_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_379.INIT_0 = 16'h0000;

ROM16 rom16_inst_380 (
    .DO(rom16_inst_380_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_380.INIT_0 = 16'h0000;

ROM16 rom16_inst_381 (
    .DO(rom16_inst_381_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_381.INIT_0 = 16'h0000;

ROM16 rom16_inst_382 (
    .DO(rom16_inst_382_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_382.INIT_0 = 16'h0000;

ROM16 rom16_inst_383 (
    .DO(rom16_inst_383_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_383.INIT_0 = 16'h0000;

ROM16 rom16_inst_384 (
    .DO(rom16_inst_384_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_384.INIT_0 = 16'h0000;

ROM16 rom16_inst_385 (
    .DO(rom16_inst_385_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_385.INIT_0 = 16'h0000;

ROM16 rom16_inst_386 (
    .DO(rom16_inst_386_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_386.INIT_0 = 16'h0000;

ROM16 rom16_inst_387 (
    .DO(rom16_inst_387_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_387.INIT_0 = 16'h0000;

ROM16 rom16_inst_388 (
    .DO(rom16_inst_388_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_388.INIT_0 = 16'h0000;

ROM16 rom16_inst_389 (
    .DO(rom16_inst_389_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_389.INIT_0 = 16'h0000;

ROM16 rom16_inst_390 (
    .DO(rom16_inst_390_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_390.INIT_0 = 16'h0000;

ROM16 rom16_inst_391 (
    .DO(rom16_inst_391_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_391.INIT_0 = 16'h0000;

ROM16 rom16_inst_392 (
    .DO(rom16_inst_392_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_392.INIT_0 = 16'h0000;

ROM16 rom16_inst_393 (
    .DO(rom16_inst_393_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_393.INIT_0 = 16'h0000;

ROM16 rom16_inst_394 (
    .DO(rom16_inst_394_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_394.INIT_0 = 16'h0000;

ROM16 rom16_inst_395 (
    .DO(rom16_inst_395_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_395.INIT_0 = 16'h0000;

ROM16 rom16_inst_396 (
    .DO(rom16_inst_396_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_396.INIT_0 = 16'h0000;

ROM16 rom16_inst_397 (
    .DO(rom16_inst_397_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_397.INIT_0 = 16'h0000;

ROM16 rom16_inst_398 (
    .DO(rom16_inst_398_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_398.INIT_0 = 16'h0000;

ROM16 rom16_inst_399 (
    .DO(rom16_inst_399_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_399.INIT_0 = 16'h0000;

ROM16 rom16_inst_400 (
    .DO(rom16_inst_400_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_400.INIT_0 = 16'h0000;

ROM16 rom16_inst_401 (
    .DO(rom16_inst_401_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_401.INIT_0 = 16'h0000;

ROM16 rom16_inst_402 (
    .DO(rom16_inst_402_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_402.INIT_0 = 16'h0000;

ROM16 rom16_inst_403 (
    .DO(rom16_inst_403_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_403.INIT_0 = 16'h0000;

ROM16 rom16_inst_404 (
    .DO(rom16_inst_404_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_404.INIT_0 = 16'h0000;

ROM16 rom16_inst_405 (
    .DO(rom16_inst_405_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_405.INIT_0 = 16'h0000;

ROM16 rom16_inst_406 (
    .DO(rom16_inst_406_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_406.INIT_0 = 16'h0000;

ROM16 rom16_inst_407 (
    .DO(rom16_inst_407_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_407.INIT_0 = 16'h0000;

ROM16 rom16_inst_408 (
    .DO(rom16_inst_408_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_408.INIT_0 = 16'h0000;

ROM16 rom16_inst_409 (
    .DO(rom16_inst_409_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_409.INIT_0 = 16'h0000;

ROM16 rom16_inst_410 (
    .DO(rom16_inst_410_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_410.INIT_0 = 16'h0000;

ROM16 rom16_inst_411 (
    .DO(rom16_inst_411_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_411.INIT_0 = 16'h0000;

ROM16 rom16_inst_412 (
    .DO(rom16_inst_412_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_412.INIT_0 = 16'h0000;

ROM16 rom16_inst_413 (
    .DO(rom16_inst_413_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_413.INIT_0 = 16'h0000;

ROM16 rom16_inst_414 (
    .DO(rom16_inst_414_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_414.INIT_0 = 16'h0000;

ROM16 rom16_inst_415 (
    .DO(rom16_inst_415_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_415.INIT_0 = 16'h0000;

ROM16 rom16_inst_416 (
    .DO(rom16_inst_416_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_416.INIT_0 = 16'h0000;

ROM16 rom16_inst_417 (
    .DO(rom16_inst_417_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_417.INIT_0 = 16'h0000;

ROM16 rom16_inst_418 (
    .DO(rom16_inst_418_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_418.INIT_0 = 16'h0000;

ROM16 rom16_inst_419 (
    .DO(rom16_inst_419_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_419.INIT_0 = 16'h0000;

ROM16 rom16_inst_420 (
    .DO(rom16_inst_420_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_420.INIT_0 = 16'h0000;

ROM16 rom16_inst_421 (
    .DO(rom16_inst_421_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_421.INIT_0 = 16'h0000;

ROM16 rom16_inst_422 (
    .DO(rom16_inst_422_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_422.INIT_0 = 16'h0000;

ROM16 rom16_inst_423 (
    .DO(rom16_inst_423_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_423.INIT_0 = 16'h0000;

ROM16 rom16_inst_424 (
    .DO(rom16_inst_424_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_424.INIT_0 = 16'h0000;

ROM16 rom16_inst_425 (
    .DO(rom16_inst_425_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_425.INIT_0 = 16'h0000;

ROM16 rom16_inst_426 (
    .DO(rom16_inst_426_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_426.INIT_0 = 16'h0000;

ROM16 rom16_inst_427 (
    .DO(rom16_inst_427_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_427.INIT_0 = 16'h0000;

ROM16 rom16_inst_428 (
    .DO(rom16_inst_428_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_428.INIT_0 = 16'h0000;

ROM16 rom16_inst_429 (
    .DO(rom16_inst_429_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_429.INIT_0 = 16'h0000;

ROM16 rom16_inst_430 (
    .DO(rom16_inst_430_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_430.INIT_0 = 16'h0000;

ROM16 rom16_inst_431 (
    .DO(rom16_inst_431_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_431.INIT_0 = 16'h0000;

ROM16 rom16_inst_432 (
    .DO(rom16_inst_432_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_432.INIT_0 = 16'h0000;

ROM16 rom16_inst_433 (
    .DO(rom16_inst_433_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_433.INIT_0 = 16'h0000;

ROM16 rom16_inst_434 (
    .DO(rom16_inst_434_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_434.INIT_0 = 16'h0000;

ROM16 rom16_inst_435 (
    .DO(rom16_inst_435_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_435.INIT_0 = 16'h0000;

ROM16 rom16_inst_436 (
    .DO(rom16_inst_436_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_436.INIT_0 = 16'h0000;

ROM16 rom16_inst_437 (
    .DO(rom16_inst_437_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_437.INIT_0 = 16'h0000;

ROM16 rom16_inst_438 (
    .DO(rom16_inst_438_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_438.INIT_0 = 16'h0000;

ROM16 rom16_inst_439 (
    .DO(rom16_inst_439_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_439.INIT_0 = 16'h0000;

ROM16 rom16_inst_440 (
    .DO(rom16_inst_440_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_440.INIT_0 = 16'h0000;

ROM16 rom16_inst_441 (
    .DO(rom16_inst_441_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_441.INIT_0 = 16'h0000;

ROM16 rom16_inst_442 (
    .DO(rom16_inst_442_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_442.INIT_0 = 16'h0000;

ROM16 rom16_inst_443 (
    .DO(rom16_inst_443_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_443.INIT_0 = 16'h0000;

ROM16 rom16_inst_444 (
    .DO(rom16_inst_444_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_444.INIT_0 = 16'h0000;

ROM16 rom16_inst_445 (
    .DO(rom16_inst_445_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_445.INIT_0 = 16'h0000;

ROM16 rom16_inst_446 (
    .DO(rom16_inst_446_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_446.INIT_0 = 16'h0000;

ROM16 rom16_inst_447 (
    .DO(rom16_inst_447_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_447.INIT_0 = 16'h0000;

ROM16 rom16_inst_448 (
    .DO(rom16_inst_448_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_448.INIT_0 = 16'h0000;

ROM16 rom16_inst_449 (
    .DO(rom16_inst_449_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_449.INIT_0 = 16'h0000;

ROM16 rom16_inst_450 (
    .DO(rom16_inst_450_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_450.INIT_0 = 16'h0000;

ROM16 rom16_inst_451 (
    .DO(rom16_inst_451_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_451.INIT_0 = 16'h0000;

ROM16 rom16_inst_452 (
    .DO(rom16_inst_452_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_452.INIT_0 = 16'h0000;

ROM16 rom16_inst_453 (
    .DO(rom16_inst_453_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_453.INIT_0 = 16'h0000;

ROM16 rom16_inst_454 (
    .DO(rom16_inst_454_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_454.INIT_0 = 16'h0000;

ROM16 rom16_inst_455 (
    .DO(rom16_inst_455_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_455.INIT_0 = 16'h0000;

ROM16 rom16_inst_456 (
    .DO(rom16_inst_456_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_456.INIT_0 = 16'h0000;

ROM16 rom16_inst_457 (
    .DO(rom16_inst_457_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_457.INIT_0 = 16'h0000;

ROM16 rom16_inst_458 (
    .DO(rom16_inst_458_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_458.INIT_0 = 16'h0000;

ROM16 rom16_inst_459 (
    .DO(rom16_inst_459_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_459.INIT_0 = 16'h0000;

ROM16 rom16_inst_460 (
    .DO(rom16_inst_460_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_460.INIT_0 = 16'h0000;

ROM16 rom16_inst_461 (
    .DO(rom16_inst_461_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_461.INIT_0 = 16'h0000;

ROM16 rom16_inst_462 (
    .DO(rom16_inst_462_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_462.INIT_0 = 16'h0000;

ROM16 rom16_inst_463 (
    .DO(rom16_inst_463_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_463.INIT_0 = 16'h0000;

ROM16 rom16_inst_464 (
    .DO(rom16_inst_464_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_464.INIT_0 = 16'h0000;

ROM16 rom16_inst_465 (
    .DO(rom16_inst_465_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_465.INIT_0 = 16'h0000;

ROM16 rom16_inst_466 (
    .DO(rom16_inst_466_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_466.INIT_0 = 16'h0000;

ROM16 rom16_inst_467 (
    .DO(rom16_inst_467_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_467.INIT_0 = 16'h0000;

ROM16 rom16_inst_468 (
    .DO(rom16_inst_468_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_468.INIT_0 = 16'h0000;

ROM16 rom16_inst_469 (
    .DO(rom16_inst_469_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_469.INIT_0 = 16'h0000;

ROM16 rom16_inst_470 (
    .DO(rom16_inst_470_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_470.INIT_0 = 16'h0000;

ROM16 rom16_inst_471 (
    .DO(rom16_inst_471_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_471.INIT_0 = 16'h0000;

ROM16 rom16_inst_472 (
    .DO(rom16_inst_472_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_472.INIT_0 = 16'h0000;

ROM16 rom16_inst_473 (
    .DO(rom16_inst_473_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_473.INIT_0 = 16'h0000;

ROM16 rom16_inst_474 (
    .DO(rom16_inst_474_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_474.INIT_0 = 16'h0000;

ROM16 rom16_inst_475 (
    .DO(rom16_inst_475_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_475.INIT_0 = 16'h0000;

ROM16 rom16_inst_476 (
    .DO(rom16_inst_476_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_476.INIT_0 = 16'h0000;

ROM16 rom16_inst_477 (
    .DO(rom16_inst_477_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_477.INIT_0 = 16'h0000;

ROM16 rom16_inst_478 (
    .DO(rom16_inst_478_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_478.INIT_0 = 16'h0000;

ROM16 rom16_inst_479 (
    .DO(rom16_inst_479_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_479.INIT_0 = 16'h0000;

ROM16 rom16_inst_480 (
    .DO(rom16_inst_480_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_480.INIT_0 = 16'h0000;

ROM16 rom16_inst_481 (
    .DO(rom16_inst_481_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_481.INIT_0 = 16'h0000;

ROM16 rom16_inst_482 (
    .DO(rom16_inst_482_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_482.INIT_0 = 16'h0000;

ROM16 rom16_inst_483 (
    .DO(rom16_inst_483_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_483.INIT_0 = 16'h0000;

ROM16 rom16_inst_484 (
    .DO(rom16_inst_484_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_484.INIT_0 = 16'h0000;

ROM16 rom16_inst_485 (
    .DO(rom16_inst_485_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_485.INIT_0 = 16'h0000;

ROM16 rom16_inst_486 (
    .DO(rom16_inst_486_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_486.INIT_0 = 16'h0000;

ROM16 rom16_inst_487 (
    .DO(rom16_inst_487_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_487.INIT_0 = 16'h0000;

ROM16 rom16_inst_488 (
    .DO(rom16_inst_488_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_488.INIT_0 = 16'h0000;

ROM16 rom16_inst_489 (
    .DO(rom16_inst_489_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_489.INIT_0 = 16'h0000;

ROM16 rom16_inst_490 (
    .DO(rom16_inst_490_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_490.INIT_0 = 16'h0000;

ROM16 rom16_inst_491 (
    .DO(rom16_inst_491_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_491.INIT_0 = 16'h0000;

ROM16 rom16_inst_492 (
    .DO(rom16_inst_492_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_492.INIT_0 = 16'h0000;

ROM16 rom16_inst_493 (
    .DO(rom16_inst_493_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_493.INIT_0 = 16'h0000;

ROM16 rom16_inst_494 (
    .DO(rom16_inst_494_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_494.INIT_0 = 16'h0000;

ROM16 rom16_inst_495 (
    .DO(rom16_inst_495_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_495.INIT_0 = 16'h0000;

ROM16 rom16_inst_496 (
    .DO(rom16_inst_496_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_496.INIT_0 = 16'h0000;

ROM16 rom16_inst_497 (
    .DO(rom16_inst_497_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_497.INIT_0 = 16'h0000;

ROM16 rom16_inst_498 (
    .DO(rom16_inst_498_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_498.INIT_0 = 16'h0000;

ROM16 rom16_inst_499 (
    .DO(rom16_inst_499_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_499.INIT_0 = 16'h0000;

ROM16 rom16_inst_500 (
    .DO(rom16_inst_500_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_500.INIT_0 = 16'h0000;

ROM16 rom16_inst_501 (
    .DO(rom16_inst_501_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_501.INIT_0 = 16'h0000;

ROM16 rom16_inst_502 (
    .DO(rom16_inst_502_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_502.INIT_0 = 16'h0000;

ROM16 rom16_inst_503 (
    .DO(rom16_inst_503_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_503.INIT_0 = 16'h0000;

ROM16 rom16_inst_504 (
    .DO(rom16_inst_504_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_504.INIT_0 = 16'h0000;

ROM16 rom16_inst_505 (
    .DO(rom16_inst_505_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_505.INIT_0 = 16'h0000;

ROM16 rom16_inst_506 (
    .DO(rom16_inst_506_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_506.INIT_0 = 16'h0000;

ROM16 rom16_inst_507 (
    .DO(rom16_inst_507_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_507.INIT_0 = 16'h0000;

ROM16 rom16_inst_508 (
    .DO(rom16_inst_508_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_508.INIT_0 = 16'h0000;

ROM16 rom16_inst_509 (
    .DO(rom16_inst_509_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_509.INIT_0 = 16'h0000;

ROM16 rom16_inst_510 (
    .DO(rom16_inst_510_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_510.INIT_0 = 16'h0000;

ROM16 rom16_inst_511 (
    .DO(rom16_inst_511_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_511.INIT_0 = 16'h0000;

ROM16 rom16_inst_512 (
    .DO(rom16_inst_512_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_512.INIT_0 = 16'h0000;

ROM16 rom16_inst_513 (
    .DO(rom16_inst_513_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_513.INIT_0 = 16'h0000;

ROM16 rom16_inst_514 (
    .DO(rom16_inst_514_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_514.INIT_0 = 16'h0000;

ROM16 rom16_inst_515 (
    .DO(rom16_inst_515_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_515.INIT_0 = 16'h0000;

ROM16 rom16_inst_516 (
    .DO(rom16_inst_516_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_516.INIT_0 = 16'h0000;

ROM16 rom16_inst_517 (
    .DO(rom16_inst_517_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_517.INIT_0 = 16'h0000;

ROM16 rom16_inst_518 (
    .DO(rom16_inst_518_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_518.INIT_0 = 16'h0000;

ROM16 rom16_inst_519 (
    .DO(rom16_inst_519_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_519.INIT_0 = 16'h0000;

ROM16 rom16_inst_520 (
    .DO(rom16_inst_520_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_520.INIT_0 = 16'h0000;

ROM16 rom16_inst_521 (
    .DO(rom16_inst_521_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_521.INIT_0 = 16'h0000;

ROM16 rom16_inst_522 (
    .DO(rom16_inst_522_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_522.INIT_0 = 16'h0000;

ROM16 rom16_inst_523 (
    .DO(rom16_inst_523_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_523.INIT_0 = 16'h0000;

ROM16 rom16_inst_524 (
    .DO(rom16_inst_524_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_524.INIT_0 = 16'h0000;

ROM16 rom16_inst_525 (
    .DO(rom16_inst_525_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_525.INIT_0 = 16'h0000;

ROM16 rom16_inst_526 (
    .DO(rom16_inst_526_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_526.INIT_0 = 16'h0000;

ROM16 rom16_inst_527 (
    .DO(rom16_inst_527_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_527.INIT_0 = 16'h0000;

ROM16 rom16_inst_528 (
    .DO(rom16_inst_528_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_528.INIT_0 = 16'h0000;

ROM16 rom16_inst_529 (
    .DO(rom16_inst_529_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_529.INIT_0 = 16'h0000;

ROM16 rom16_inst_530 (
    .DO(rom16_inst_530_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_530.INIT_0 = 16'h0000;

ROM16 rom16_inst_531 (
    .DO(rom16_inst_531_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_531.INIT_0 = 16'h0000;

ROM16 rom16_inst_532 (
    .DO(rom16_inst_532_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_532.INIT_0 = 16'h0000;

ROM16 rom16_inst_533 (
    .DO(rom16_inst_533_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_533.INIT_0 = 16'h0000;

ROM16 rom16_inst_534 (
    .DO(rom16_inst_534_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_534.INIT_0 = 16'h0000;

ROM16 rom16_inst_535 (
    .DO(rom16_inst_535_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_535.INIT_0 = 16'h0000;

ROM16 rom16_inst_536 (
    .DO(rom16_inst_536_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_536.INIT_0 = 16'h0000;

ROM16 rom16_inst_537 (
    .DO(rom16_inst_537_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_537.INIT_0 = 16'h0000;

ROM16 rom16_inst_538 (
    .DO(rom16_inst_538_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_538.INIT_0 = 16'h0000;

ROM16 rom16_inst_539 (
    .DO(rom16_inst_539_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_539.INIT_0 = 16'h0000;

ROM16 rom16_inst_540 (
    .DO(rom16_inst_540_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_540.INIT_0 = 16'h0000;

ROM16 rom16_inst_541 (
    .DO(rom16_inst_541_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_541.INIT_0 = 16'h0000;

ROM16 rom16_inst_542 (
    .DO(rom16_inst_542_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_542.INIT_0 = 16'h0000;

ROM16 rom16_inst_543 (
    .DO(rom16_inst_543_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_543.INIT_0 = 16'h0000;

ROM16 rom16_inst_544 (
    .DO(rom16_inst_544_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_544.INIT_0 = 16'h0000;

ROM16 rom16_inst_545 (
    .DO(rom16_inst_545_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_545.INIT_0 = 16'h0000;

ROM16 rom16_inst_546 (
    .DO(rom16_inst_546_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_546.INIT_0 = 16'h0000;

ROM16 rom16_inst_547 (
    .DO(rom16_inst_547_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_547.INIT_0 = 16'h0000;

ROM16 rom16_inst_548 (
    .DO(rom16_inst_548_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_548.INIT_0 = 16'h0000;

ROM16 rom16_inst_549 (
    .DO(rom16_inst_549_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_549.INIT_0 = 16'h0000;

ROM16 rom16_inst_550 (
    .DO(rom16_inst_550_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_550.INIT_0 = 16'h0000;

ROM16 rom16_inst_551 (
    .DO(rom16_inst_551_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_551.INIT_0 = 16'h0000;

ROM16 rom16_inst_552 (
    .DO(rom16_inst_552_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_552.INIT_0 = 16'h0000;

ROM16 rom16_inst_553 (
    .DO(rom16_inst_553_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_553.INIT_0 = 16'h0000;

ROM16 rom16_inst_554 (
    .DO(rom16_inst_554_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_554.INIT_0 = 16'h0000;

ROM16 rom16_inst_555 (
    .DO(rom16_inst_555_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_555.INIT_0 = 16'h0000;

ROM16 rom16_inst_556 (
    .DO(rom16_inst_556_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_556.INIT_0 = 16'h0000;

ROM16 rom16_inst_557 (
    .DO(rom16_inst_557_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_557.INIT_0 = 16'h0000;

ROM16 rom16_inst_558 (
    .DO(rom16_inst_558_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_558.INIT_0 = 16'h0000;

ROM16 rom16_inst_559 (
    .DO(rom16_inst_559_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_559.INIT_0 = 16'h0000;

ROM16 rom16_inst_560 (
    .DO(rom16_inst_560_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_560.INIT_0 = 16'h0000;

ROM16 rom16_inst_561 (
    .DO(rom16_inst_561_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_561.INIT_0 = 16'h0000;

ROM16 rom16_inst_562 (
    .DO(rom16_inst_562_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_562.INIT_0 = 16'h0000;

ROM16 rom16_inst_563 (
    .DO(rom16_inst_563_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_563.INIT_0 = 16'h0000;

ROM16 rom16_inst_564 (
    .DO(rom16_inst_564_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_564.INIT_0 = 16'h0000;

ROM16 rom16_inst_565 (
    .DO(rom16_inst_565_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_565.INIT_0 = 16'h0000;

ROM16 rom16_inst_566 (
    .DO(rom16_inst_566_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_566.INIT_0 = 16'h0000;

ROM16 rom16_inst_567 (
    .DO(rom16_inst_567_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_567.INIT_0 = 16'h0000;

ROM16 rom16_inst_568 (
    .DO(rom16_inst_568_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_568.INIT_0 = 16'h0000;

ROM16 rom16_inst_569 (
    .DO(rom16_inst_569_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_569.INIT_0 = 16'h0000;

ROM16 rom16_inst_570 (
    .DO(rom16_inst_570_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_570.INIT_0 = 16'h0000;

ROM16 rom16_inst_571 (
    .DO(rom16_inst_571_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_571.INIT_0 = 16'h0000;

ROM16 rom16_inst_572 (
    .DO(rom16_inst_572_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_572.INIT_0 = 16'h0000;

ROM16 rom16_inst_573 (
    .DO(rom16_inst_573_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_573.INIT_0 = 16'h0000;

ROM16 rom16_inst_574 (
    .DO(rom16_inst_574_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_574.INIT_0 = 16'h0000;

ROM16 rom16_inst_575 (
    .DO(rom16_inst_575_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_575.INIT_0 = 16'h0000;

ROM16 rom16_inst_576 (
    .DO(rom16_inst_576_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_576.INIT_0 = 16'h0000;

ROM16 rom16_inst_577 (
    .DO(rom16_inst_577_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_577.INIT_0 = 16'h0000;

ROM16 rom16_inst_578 (
    .DO(rom16_inst_578_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_578.INIT_0 = 16'h0000;

ROM16 rom16_inst_579 (
    .DO(rom16_inst_579_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_579.INIT_0 = 16'h0000;

ROM16 rom16_inst_580 (
    .DO(rom16_inst_580_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_580.INIT_0 = 16'h0000;

ROM16 rom16_inst_581 (
    .DO(rom16_inst_581_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_581.INIT_0 = 16'h0000;

ROM16 rom16_inst_582 (
    .DO(rom16_inst_582_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_582.INIT_0 = 16'h0000;

ROM16 rom16_inst_583 (
    .DO(rom16_inst_583_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_583.INIT_0 = 16'h0000;

ROM16 rom16_inst_584 (
    .DO(rom16_inst_584_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_584.INIT_0 = 16'h0000;

ROM16 rom16_inst_585 (
    .DO(rom16_inst_585_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_585.INIT_0 = 16'h0000;

ROM16 rom16_inst_586 (
    .DO(rom16_inst_586_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_586.INIT_0 = 16'h0000;

ROM16 rom16_inst_587 (
    .DO(rom16_inst_587_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_587.INIT_0 = 16'h0000;

ROM16 rom16_inst_588 (
    .DO(rom16_inst_588_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_588.INIT_0 = 16'h0000;

ROM16 rom16_inst_589 (
    .DO(rom16_inst_589_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_589.INIT_0 = 16'h0000;

ROM16 rom16_inst_590 (
    .DO(rom16_inst_590_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_590.INIT_0 = 16'h0000;

ROM16 rom16_inst_591 (
    .DO(rom16_inst_591_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_591.INIT_0 = 16'h0000;

ROM16 rom16_inst_592 (
    .DO(rom16_inst_592_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_592.INIT_0 = 16'h0000;

ROM16 rom16_inst_593 (
    .DO(rom16_inst_593_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_593.INIT_0 = 16'h0000;

ROM16 rom16_inst_594 (
    .DO(rom16_inst_594_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_594.INIT_0 = 16'h0000;

ROM16 rom16_inst_595 (
    .DO(rom16_inst_595_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_595.INIT_0 = 16'h0000;

ROM16 rom16_inst_596 (
    .DO(rom16_inst_596_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_596.INIT_0 = 16'h0000;

ROM16 rom16_inst_597 (
    .DO(rom16_inst_597_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_597.INIT_0 = 16'h0000;

ROM16 rom16_inst_598 (
    .DO(rom16_inst_598_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_598.INIT_0 = 16'h0000;

ROM16 rom16_inst_599 (
    .DO(rom16_inst_599_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_599.INIT_0 = 16'h0000;

ROM16 rom16_inst_600 (
    .DO(rom16_inst_600_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_600.INIT_0 = 16'h0000;

ROM16 rom16_inst_601 (
    .DO(rom16_inst_601_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_601.INIT_0 = 16'h0000;

ROM16 rom16_inst_602 (
    .DO(rom16_inst_602_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_602.INIT_0 = 16'h0000;

ROM16 rom16_inst_603 (
    .DO(rom16_inst_603_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_603.INIT_0 = 16'h0000;

ROM16 rom16_inst_604 (
    .DO(rom16_inst_604_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_604.INIT_0 = 16'h0000;

ROM16 rom16_inst_605 (
    .DO(rom16_inst_605_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_605.INIT_0 = 16'h0000;

ROM16 rom16_inst_606 (
    .DO(rom16_inst_606_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_606.INIT_0 = 16'h0000;

ROM16 rom16_inst_607 (
    .DO(rom16_inst_607_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_607.INIT_0 = 16'h0000;

ROM16 rom16_inst_608 (
    .DO(rom16_inst_608_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_608.INIT_0 = 16'h0000;

ROM16 rom16_inst_609 (
    .DO(rom16_inst_609_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_609.INIT_0 = 16'h0000;

ROM16 rom16_inst_610 (
    .DO(rom16_inst_610_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_610.INIT_0 = 16'h0000;

ROM16 rom16_inst_611 (
    .DO(rom16_inst_611_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_611.INIT_0 = 16'h0000;

ROM16 rom16_inst_612 (
    .DO(rom16_inst_612_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_612.INIT_0 = 16'h0000;

ROM16 rom16_inst_613 (
    .DO(rom16_inst_613_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_613.INIT_0 = 16'h0000;

ROM16 rom16_inst_614 (
    .DO(rom16_inst_614_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_614.INIT_0 = 16'h0000;

ROM16 rom16_inst_615 (
    .DO(rom16_inst_615_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_615.INIT_0 = 16'h0000;

ROM16 rom16_inst_616 (
    .DO(rom16_inst_616_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_616.INIT_0 = 16'h0000;

ROM16 rom16_inst_617 (
    .DO(rom16_inst_617_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_617.INIT_0 = 16'h0000;

ROM16 rom16_inst_618 (
    .DO(rom16_inst_618_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_618.INIT_0 = 16'h0000;

ROM16 rom16_inst_619 (
    .DO(rom16_inst_619_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_619.INIT_0 = 16'h0000;

ROM16 rom16_inst_620 (
    .DO(rom16_inst_620_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_620.INIT_0 = 16'h0000;

ROM16 rom16_inst_621 (
    .DO(rom16_inst_621_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_621.INIT_0 = 16'h0000;

ROM16 rom16_inst_622 (
    .DO(rom16_inst_622_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_622.INIT_0 = 16'h0000;

ROM16 rom16_inst_623 (
    .DO(rom16_inst_623_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_623.INIT_0 = 16'h0000;

ROM16 rom16_inst_624 (
    .DO(rom16_inst_624_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_624.INIT_0 = 16'h0000;

ROM16 rom16_inst_625 (
    .DO(rom16_inst_625_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_625.INIT_0 = 16'h0000;

ROM16 rom16_inst_626 (
    .DO(rom16_inst_626_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_626.INIT_0 = 16'h0000;

ROM16 rom16_inst_627 (
    .DO(rom16_inst_627_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_627.INIT_0 = 16'h0000;

ROM16 rom16_inst_628 (
    .DO(rom16_inst_628_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_628.INIT_0 = 16'h0000;

ROM16 rom16_inst_629 (
    .DO(rom16_inst_629_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_629.INIT_0 = 16'h0000;

ROM16 rom16_inst_630 (
    .DO(rom16_inst_630_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_630.INIT_0 = 16'h0000;

ROM16 rom16_inst_631 (
    .DO(rom16_inst_631_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_631.INIT_0 = 16'h0000;

ROM16 rom16_inst_632 (
    .DO(rom16_inst_632_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_632.INIT_0 = 16'h0000;

ROM16 rom16_inst_633 (
    .DO(rom16_inst_633_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_633.INIT_0 = 16'h0000;

ROM16 rom16_inst_634 (
    .DO(rom16_inst_634_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_634.INIT_0 = 16'h0000;

ROM16 rom16_inst_635 (
    .DO(rom16_inst_635_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_635.INIT_0 = 16'h0000;

ROM16 rom16_inst_636 (
    .DO(rom16_inst_636_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_636.INIT_0 = 16'h0000;

ROM16 rom16_inst_637 (
    .DO(rom16_inst_637_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_637.INIT_0 = 16'h0000;

ROM16 rom16_inst_638 (
    .DO(rom16_inst_638_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_638.INIT_0 = 16'h0000;

ROM16 rom16_inst_639 (
    .DO(rom16_inst_639_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_639.INIT_0 = 16'h0000;

ROM16 rom16_inst_640 (
    .DO(rom16_inst_640_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_640.INIT_0 = 16'h0000;

ROM16 rom16_inst_641 (
    .DO(rom16_inst_641_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_641.INIT_0 = 16'h0000;

ROM16 rom16_inst_642 (
    .DO(rom16_inst_642_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_642.INIT_0 = 16'h0000;

ROM16 rom16_inst_643 (
    .DO(rom16_inst_643_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_643.INIT_0 = 16'h0000;

ROM16 rom16_inst_644 (
    .DO(rom16_inst_644_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_644.INIT_0 = 16'h0000;

ROM16 rom16_inst_645 (
    .DO(rom16_inst_645_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_645.INIT_0 = 16'h0000;

ROM16 rom16_inst_646 (
    .DO(rom16_inst_646_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_646.INIT_0 = 16'h0000;

ROM16 rom16_inst_647 (
    .DO(rom16_inst_647_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_647.INIT_0 = 16'h0000;

ROM16 rom16_inst_648 (
    .DO(rom16_inst_648_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_648.INIT_0 = 16'h0000;

ROM16 rom16_inst_649 (
    .DO(rom16_inst_649_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_649.INIT_0 = 16'h0000;

ROM16 rom16_inst_650 (
    .DO(rom16_inst_650_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_650.INIT_0 = 16'h0000;

ROM16 rom16_inst_651 (
    .DO(rom16_inst_651_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_651.INIT_0 = 16'h0000;

ROM16 rom16_inst_652 (
    .DO(rom16_inst_652_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_652.INIT_0 = 16'h0000;

ROM16 rom16_inst_653 (
    .DO(rom16_inst_653_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_653.INIT_0 = 16'h0000;

ROM16 rom16_inst_654 (
    .DO(rom16_inst_654_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_654.INIT_0 = 16'h0000;

ROM16 rom16_inst_655 (
    .DO(rom16_inst_655_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_655.INIT_0 = 16'h0000;

ROM16 rom16_inst_656 (
    .DO(rom16_inst_656_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_656.INIT_0 = 16'h0000;

ROM16 rom16_inst_657 (
    .DO(rom16_inst_657_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_657.INIT_0 = 16'h0000;

ROM16 rom16_inst_658 (
    .DO(rom16_inst_658_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_658.INIT_0 = 16'h0000;

ROM16 rom16_inst_659 (
    .DO(rom16_inst_659_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_659.INIT_0 = 16'h0000;

ROM16 rom16_inst_660 (
    .DO(rom16_inst_660_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_660.INIT_0 = 16'h0000;

ROM16 rom16_inst_661 (
    .DO(rom16_inst_661_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_661.INIT_0 = 16'h0000;

ROM16 rom16_inst_662 (
    .DO(rom16_inst_662_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_662.INIT_0 = 16'h0000;

ROM16 rom16_inst_663 (
    .DO(rom16_inst_663_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_663.INIT_0 = 16'h0000;

ROM16 rom16_inst_664 (
    .DO(rom16_inst_664_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_664.INIT_0 = 16'h0000;

ROM16 rom16_inst_665 (
    .DO(rom16_inst_665_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_665.INIT_0 = 16'h0000;

ROM16 rom16_inst_666 (
    .DO(rom16_inst_666_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_666.INIT_0 = 16'h0000;

ROM16 rom16_inst_667 (
    .DO(rom16_inst_667_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_667.INIT_0 = 16'h0000;

ROM16 rom16_inst_668 (
    .DO(rom16_inst_668_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_668.INIT_0 = 16'h0000;

ROM16 rom16_inst_669 (
    .DO(rom16_inst_669_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_669.INIT_0 = 16'h0000;

ROM16 rom16_inst_670 (
    .DO(rom16_inst_670_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_670.INIT_0 = 16'h0000;

ROM16 rom16_inst_671 (
    .DO(rom16_inst_671_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_671.INIT_0 = 16'h0000;

ROM16 rom16_inst_672 (
    .DO(rom16_inst_672_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_672.INIT_0 = 16'h0000;

ROM16 rom16_inst_673 (
    .DO(rom16_inst_673_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_673.INIT_0 = 16'h0000;

ROM16 rom16_inst_674 (
    .DO(rom16_inst_674_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_674.INIT_0 = 16'h0000;

ROM16 rom16_inst_675 (
    .DO(rom16_inst_675_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_675.INIT_0 = 16'h0000;

ROM16 rom16_inst_676 (
    .DO(rom16_inst_676_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_676.INIT_0 = 16'h0000;

ROM16 rom16_inst_677 (
    .DO(rom16_inst_677_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_677.INIT_0 = 16'h0000;

ROM16 rom16_inst_678 (
    .DO(rom16_inst_678_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_678.INIT_0 = 16'h0000;

ROM16 rom16_inst_679 (
    .DO(rom16_inst_679_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_679.INIT_0 = 16'h0000;

ROM16 rom16_inst_680 (
    .DO(rom16_inst_680_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_680.INIT_0 = 16'h0000;

ROM16 rom16_inst_681 (
    .DO(rom16_inst_681_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_681.INIT_0 = 16'h0000;

ROM16 rom16_inst_682 (
    .DO(rom16_inst_682_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_682.INIT_0 = 16'h0000;

ROM16 rom16_inst_683 (
    .DO(rom16_inst_683_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_683.INIT_0 = 16'h0000;

ROM16 rom16_inst_684 (
    .DO(rom16_inst_684_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_684.INIT_0 = 16'h0000;

ROM16 rom16_inst_685 (
    .DO(rom16_inst_685_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_685.INIT_0 = 16'h0000;

ROM16 rom16_inst_686 (
    .DO(rom16_inst_686_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_686.INIT_0 = 16'h0000;

ROM16 rom16_inst_687 (
    .DO(rom16_inst_687_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_687.INIT_0 = 16'h0000;

ROM16 rom16_inst_688 (
    .DO(rom16_inst_688_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_688.INIT_0 = 16'h0000;

ROM16 rom16_inst_689 (
    .DO(rom16_inst_689_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_689.INIT_0 = 16'h0000;

ROM16 rom16_inst_690 (
    .DO(rom16_inst_690_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_690.INIT_0 = 16'h0000;

ROM16 rom16_inst_691 (
    .DO(rom16_inst_691_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_691.INIT_0 = 16'h0000;

ROM16 rom16_inst_692 (
    .DO(rom16_inst_692_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_692.INIT_0 = 16'h0000;

ROM16 rom16_inst_693 (
    .DO(rom16_inst_693_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_693.INIT_0 = 16'h0000;

ROM16 rom16_inst_694 (
    .DO(rom16_inst_694_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_694.INIT_0 = 16'h0000;

ROM16 rom16_inst_695 (
    .DO(rom16_inst_695_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_695.INIT_0 = 16'h0000;

ROM16 rom16_inst_696 (
    .DO(rom16_inst_696_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_696.INIT_0 = 16'h0000;

ROM16 rom16_inst_697 (
    .DO(rom16_inst_697_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_697.INIT_0 = 16'h0000;

ROM16 rom16_inst_698 (
    .DO(rom16_inst_698_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_698.INIT_0 = 16'h0000;

ROM16 rom16_inst_699 (
    .DO(rom16_inst_699_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_699.INIT_0 = 16'h0000;

ROM16 rom16_inst_700 (
    .DO(rom16_inst_700_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_700.INIT_0 = 16'h0000;

ROM16 rom16_inst_701 (
    .DO(rom16_inst_701_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_701.INIT_0 = 16'h0000;

ROM16 rom16_inst_702 (
    .DO(rom16_inst_702_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_702.INIT_0 = 16'h0000;

ROM16 rom16_inst_703 (
    .DO(rom16_inst_703_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_703.INIT_0 = 16'h0000;

ROM16 rom16_inst_704 (
    .DO(rom16_inst_704_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_704.INIT_0 = 16'h0000;

ROM16 rom16_inst_705 (
    .DO(rom16_inst_705_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_705.INIT_0 = 16'h0000;

ROM16 rom16_inst_706 (
    .DO(rom16_inst_706_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_706.INIT_0 = 16'h0000;

ROM16 rom16_inst_707 (
    .DO(rom16_inst_707_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_707.INIT_0 = 16'h0000;

ROM16 rom16_inst_708 (
    .DO(rom16_inst_708_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_708.INIT_0 = 16'h0000;

ROM16 rom16_inst_709 (
    .DO(rom16_inst_709_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_709.INIT_0 = 16'h0000;

ROM16 rom16_inst_710 (
    .DO(rom16_inst_710_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_710.INIT_0 = 16'h0000;

ROM16 rom16_inst_711 (
    .DO(rom16_inst_711_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_711.INIT_0 = 16'h0000;

ROM16 rom16_inst_712 (
    .DO(rom16_inst_712_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_712.INIT_0 = 16'h0000;

ROM16 rom16_inst_713 (
    .DO(rom16_inst_713_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_713.INIT_0 = 16'h0000;

ROM16 rom16_inst_714 (
    .DO(rom16_inst_714_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_714.INIT_0 = 16'h0000;

ROM16 rom16_inst_715 (
    .DO(rom16_inst_715_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_715.INIT_0 = 16'h0000;

ROM16 rom16_inst_716 (
    .DO(rom16_inst_716_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_716.INIT_0 = 16'h0000;

ROM16 rom16_inst_717 (
    .DO(rom16_inst_717_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_717.INIT_0 = 16'h0000;

ROM16 rom16_inst_718 (
    .DO(rom16_inst_718_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_718.INIT_0 = 16'h0000;

ROM16 rom16_inst_719 (
    .DO(rom16_inst_719_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_719.INIT_0 = 16'h0000;

ROM16 rom16_inst_720 (
    .DO(rom16_inst_720_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_720.INIT_0 = 16'h0000;

ROM16 rom16_inst_721 (
    .DO(rom16_inst_721_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_721.INIT_0 = 16'h0000;

ROM16 rom16_inst_722 (
    .DO(rom16_inst_722_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_722.INIT_0 = 16'h0000;

ROM16 rom16_inst_723 (
    .DO(rom16_inst_723_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_723.INIT_0 = 16'h0000;

ROM16 rom16_inst_724 (
    .DO(rom16_inst_724_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_724.INIT_0 = 16'h0000;

ROM16 rom16_inst_725 (
    .DO(rom16_inst_725_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_725.INIT_0 = 16'h0000;

ROM16 rom16_inst_726 (
    .DO(rom16_inst_726_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_726.INIT_0 = 16'h0000;

ROM16 rom16_inst_727 (
    .DO(rom16_inst_727_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_727.INIT_0 = 16'h0000;

ROM16 rom16_inst_728 (
    .DO(rom16_inst_728_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_728.INIT_0 = 16'h0000;

ROM16 rom16_inst_729 (
    .DO(rom16_inst_729_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_729.INIT_0 = 16'h0000;

ROM16 rom16_inst_730 (
    .DO(rom16_inst_730_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_730.INIT_0 = 16'h0000;

ROM16 rom16_inst_731 (
    .DO(rom16_inst_731_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_731.INIT_0 = 16'h0000;

ROM16 rom16_inst_732 (
    .DO(rom16_inst_732_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_732.INIT_0 = 16'h0000;

ROM16 rom16_inst_733 (
    .DO(rom16_inst_733_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_733.INIT_0 = 16'h0000;

ROM16 rom16_inst_734 (
    .DO(rom16_inst_734_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_734.INIT_0 = 16'h0000;

ROM16 rom16_inst_735 (
    .DO(rom16_inst_735_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_735.INIT_0 = 16'h0000;

ROM16 rom16_inst_736 (
    .DO(rom16_inst_736_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_736.INIT_0 = 16'h0000;

ROM16 rom16_inst_737 (
    .DO(rom16_inst_737_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_737.INIT_0 = 16'h0000;

ROM16 rom16_inst_738 (
    .DO(rom16_inst_738_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_738.INIT_0 = 16'h0000;

ROM16 rom16_inst_739 (
    .DO(rom16_inst_739_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_739.INIT_0 = 16'h0000;

ROM16 rom16_inst_740 (
    .DO(rom16_inst_740_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_740.INIT_0 = 16'h0000;

ROM16 rom16_inst_741 (
    .DO(rom16_inst_741_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_741.INIT_0 = 16'h0000;

ROM16 rom16_inst_742 (
    .DO(rom16_inst_742_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_742.INIT_0 = 16'h0000;

ROM16 rom16_inst_743 (
    .DO(rom16_inst_743_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_743.INIT_0 = 16'h0000;

ROM16 rom16_inst_744 (
    .DO(rom16_inst_744_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_744.INIT_0 = 16'h0000;

ROM16 rom16_inst_745 (
    .DO(rom16_inst_745_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_745.INIT_0 = 16'h0000;

ROM16 rom16_inst_746 (
    .DO(rom16_inst_746_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_746.INIT_0 = 16'h0000;

ROM16 rom16_inst_747 (
    .DO(rom16_inst_747_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_747.INIT_0 = 16'h0000;

ROM16 rom16_inst_748 (
    .DO(rom16_inst_748_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_748.INIT_0 = 16'h0000;

ROM16 rom16_inst_749 (
    .DO(rom16_inst_749_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_749.INIT_0 = 16'h0000;

ROM16 rom16_inst_750 (
    .DO(rom16_inst_750_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_750.INIT_0 = 16'h0000;

ROM16 rom16_inst_751 (
    .DO(rom16_inst_751_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_751.INIT_0 = 16'h0000;

ROM16 rom16_inst_752 (
    .DO(rom16_inst_752_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_752.INIT_0 = 16'h0000;

ROM16 rom16_inst_753 (
    .DO(rom16_inst_753_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_753.INIT_0 = 16'h0000;

ROM16 rom16_inst_754 (
    .DO(rom16_inst_754_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_754.INIT_0 = 16'h0000;

ROM16 rom16_inst_755 (
    .DO(rom16_inst_755_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_755.INIT_0 = 16'h0000;

ROM16 rom16_inst_756 (
    .DO(rom16_inst_756_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_756.INIT_0 = 16'h0000;

ROM16 rom16_inst_757 (
    .DO(rom16_inst_757_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_757.INIT_0 = 16'h0000;

ROM16 rom16_inst_758 (
    .DO(rom16_inst_758_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_758.INIT_0 = 16'h0000;

ROM16 rom16_inst_759 (
    .DO(rom16_inst_759_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_759.INIT_0 = 16'h0000;

ROM16 rom16_inst_760 (
    .DO(rom16_inst_760_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_760.INIT_0 = 16'h0000;

ROM16 rom16_inst_761 (
    .DO(rom16_inst_761_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_761.INIT_0 = 16'h0000;

ROM16 rom16_inst_762 (
    .DO(rom16_inst_762_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_762.INIT_0 = 16'h0000;

ROM16 rom16_inst_763 (
    .DO(rom16_inst_763_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_763.INIT_0 = 16'h0000;

ROM16 rom16_inst_764 (
    .DO(rom16_inst_764_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_764.INIT_0 = 16'h0000;

ROM16 rom16_inst_765 (
    .DO(rom16_inst_765_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_765.INIT_0 = 16'h0000;

ROM16 rom16_inst_766 (
    .DO(rom16_inst_766_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_766.INIT_0 = 16'h0000;

ROM16 rom16_inst_767 (
    .DO(rom16_inst_767_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_767.INIT_0 = 16'h0000;

ROM16 rom16_inst_768 (
    .DO(rom16_inst_768_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_768.INIT_0 = 16'h0000;

ROM16 rom16_inst_769 (
    .DO(rom16_inst_769_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_769.INIT_0 = 16'h0000;

ROM16 rom16_inst_770 (
    .DO(rom16_inst_770_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_770.INIT_0 = 16'h0000;

ROM16 rom16_inst_771 (
    .DO(rom16_inst_771_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_771.INIT_0 = 16'h0000;

ROM16 rom16_inst_772 (
    .DO(rom16_inst_772_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_772.INIT_0 = 16'h0000;

ROM16 rom16_inst_773 (
    .DO(rom16_inst_773_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_773.INIT_0 = 16'h0000;

ROM16 rom16_inst_774 (
    .DO(rom16_inst_774_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_774.INIT_0 = 16'h0000;

ROM16 rom16_inst_775 (
    .DO(rom16_inst_775_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_775.INIT_0 = 16'h0000;

ROM16 rom16_inst_776 (
    .DO(rom16_inst_776_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_776.INIT_0 = 16'h0000;

ROM16 rom16_inst_777 (
    .DO(rom16_inst_777_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_777.INIT_0 = 16'h0000;

ROM16 rom16_inst_778 (
    .DO(rom16_inst_778_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_778.INIT_0 = 16'h0000;

ROM16 rom16_inst_779 (
    .DO(rom16_inst_779_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_779.INIT_0 = 16'h0000;

ROM16 rom16_inst_780 (
    .DO(rom16_inst_780_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_780.INIT_0 = 16'h0000;

ROM16 rom16_inst_781 (
    .DO(rom16_inst_781_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_781.INIT_0 = 16'h0000;

ROM16 rom16_inst_782 (
    .DO(rom16_inst_782_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_782.INIT_0 = 16'h0000;

ROM16 rom16_inst_783 (
    .DO(rom16_inst_783_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_783.INIT_0 = 16'h0000;

ROM16 rom16_inst_784 (
    .DO(rom16_inst_784_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_784.INIT_0 = 16'h0000;

ROM16 rom16_inst_785 (
    .DO(rom16_inst_785_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_785.INIT_0 = 16'h0000;

ROM16 rom16_inst_786 (
    .DO(rom16_inst_786_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_786.INIT_0 = 16'h0000;

ROM16 rom16_inst_787 (
    .DO(rom16_inst_787_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_787.INIT_0 = 16'h0000;

ROM16 rom16_inst_788 (
    .DO(rom16_inst_788_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_788.INIT_0 = 16'h0000;

ROM16 rom16_inst_789 (
    .DO(rom16_inst_789_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_789.INIT_0 = 16'h0000;

ROM16 rom16_inst_790 (
    .DO(rom16_inst_790_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_790.INIT_0 = 16'h0000;

ROM16 rom16_inst_791 (
    .DO(rom16_inst_791_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_791.INIT_0 = 16'h0000;

ROM16 rom16_inst_792 (
    .DO(rom16_inst_792_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_792.INIT_0 = 16'h0000;

ROM16 rom16_inst_793 (
    .DO(rom16_inst_793_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_793.INIT_0 = 16'h0000;

ROM16 rom16_inst_794 (
    .DO(rom16_inst_794_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_794.INIT_0 = 16'h0000;

ROM16 rom16_inst_795 (
    .DO(rom16_inst_795_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_795.INIT_0 = 16'h0000;

ROM16 rom16_inst_796 (
    .DO(rom16_inst_796_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_796.INIT_0 = 16'h0000;

ROM16 rom16_inst_797 (
    .DO(rom16_inst_797_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_797.INIT_0 = 16'h0000;

ROM16 rom16_inst_798 (
    .DO(rom16_inst_798_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_798.INIT_0 = 16'h0000;

ROM16 rom16_inst_799 (
    .DO(rom16_inst_799_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_799.INIT_0 = 16'h0000;

ROM16 rom16_inst_800 (
    .DO(rom16_inst_800_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_800.INIT_0 = 16'h0000;

ROM16 rom16_inst_801 (
    .DO(rom16_inst_801_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_801.INIT_0 = 16'h0000;

ROM16 rom16_inst_802 (
    .DO(rom16_inst_802_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_802.INIT_0 = 16'h0000;

ROM16 rom16_inst_803 (
    .DO(rom16_inst_803_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_803.INIT_0 = 16'h0000;

ROM16 rom16_inst_804 (
    .DO(rom16_inst_804_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_804.INIT_0 = 16'h0000;

ROM16 rom16_inst_805 (
    .DO(rom16_inst_805_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_805.INIT_0 = 16'h0000;

ROM16 rom16_inst_806 (
    .DO(rom16_inst_806_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_806.INIT_0 = 16'h0000;

ROM16 rom16_inst_807 (
    .DO(rom16_inst_807_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_807.INIT_0 = 16'h0000;

ROM16 rom16_inst_808 (
    .DO(rom16_inst_808_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_808.INIT_0 = 16'h0000;

ROM16 rom16_inst_809 (
    .DO(rom16_inst_809_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_809.INIT_0 = 16'h0000;

ROM16 rom16_inst_810 (
    .DO(rom16_inst_810_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_810.INIT_0 = 16'h0000;

ROM16 rom16_inst_811 (
    .DO(rom16_inst_811_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_811.INIT_0 = 16'h0000;

ROM16 rom16_inst_812 (
    .DO(rom16_inst_812_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_812.INIT_0 = 16'h0000;

ROM16 rom16_inst_813 (
    .DO(rom16_inst_813_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_813.INIT_0 = 16'h0000;

ROM16 rom16_inst_814 (
    .DO(rom16_inst_814_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_814.INIT_0 = 16'h0000;

ROM16 rom16_inst_815 (
    .DO(rom16_inst_815_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_815.INIT_0 = 16'h0000;

ROM16 rom16_inst_816 (
    .DO(rom16_inst_816_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_816.INIT_0 = 16'h0000;

ROM16 rom16_inst_817 (
    .DO(rom16_inst_817_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_817.INIT_0 = 16'h0000;

ROM16 rom16_inst_818 (
    .DO(rom16_inst_818_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_818.INIT_0 = 16'h0000;

ROM16 rom16_inst_819 (
    .DO(rom16_inst_819_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_819.INIT_0 = 16'h0000;

ROM16 rom16_inst_820 (
    .DO(rom16_inst_820_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_820.INIT_0 = 16'h0000;

ROM16 rom16_inst_821 (
    .DO(rom16_inst_821_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_821.INIT_0 = 16'h0000;

ROM16 rom16_inst_822 (
    .DO(rom16_inst_822_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_822.INIT_0 = 16'h0000;

ROM16 rom16_inst_823 (
    .DO(rom16_inst_823_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_823.INIT_0 = 16'h0000;

ROM16 rom16_inst_824 (
    .DO(rom16_inst_824_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_824.INIT_0 = 16'h0000;

ROM16 rom16_inst_825 (
    .DO(rom16_inst_825_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_825.INIT_0 = 16'h0000;

ROM16 rom16_inst_826 (
    .DO(rom16_inst_826_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_826.INIT_0 = 16'h0000;

ROM16 rom16_inst_827 (
    .DO(rom16_inst_827_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_827.INIT_0 = 16'h0000;

ROM16 rom16_inst_828 (
    .DO(rom16_inst_828_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_828.INIT_0 = 16'h0000;

ROM16 rom16_inst_829 (
    .DO(rom16_inst_829_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_829.INIT_0 = 16'h0000;

ROM16 rom16_inst_830 (
    .DO(rom16_inst_830_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_830.INIT_0 = 16'h0000;

ROM16 rom16_inst_831 (
    .DO(rom16_inst_831_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_831.INIT_0 = 16'h0000;

ROM16 rom16_inst_832 (
    .DO(rom16_inst_832_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_832.INIT_0 = 16'h0000;

ROM16 rom16_inst_833 (
    .DO(rom16_inst_833_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_833.INIT_0 = 16'h0000;

ROM16 rom16_inst_834 (
    .DO(rom16_inst_834_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_834.INIT_0 = 16'h0000;

ROM16 rom16_inst_835 (
    .DO(rom16_inst_835_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_835.INIT_0 = 16'h0000;

ROM16 rom16_inst_836 (
    .DO(rom16_inst_836_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_836.INIT_0 = 16'h0000;

ROM16 rom16_inst_837 (
    .DO(rom16_inst_837_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_837.INIT_0 = 16'h0000;

ROM16 rom16_inst_838 (
    .DO(rom16_inst_838_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_838.INIT_0 = 16'h0000;

ROM16 rom16_inst_839 (
    .DO(rom16_inst_839_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_839.INIT_0 = 16'h0000;

ROM16 rom16_inst_840 (
    .DO(rom16_inst_840_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_840.INIT_0 = 16'h0000;

ROM16 rom16_inst_841 (
    .DO(rom16_inst_841_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_841.INIT_0 = 16'h0000;

ROM16 rom16_inst_842 (
    .DO(rom16_inst_842_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_842.INIT_0 = 16'h0000;

ROM16 rom16_inst_843 (
    .DO(rom16_inst_843_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_843.INIT_0 = 16'h0000;

ROM16 rom16_inst_844 (
    .DO(rom16_inst_844_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_844.INIT_0 = 16'h0000;

ROM16 rom16_inst_845 (
    .DO(rom16_inst_845_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_845.INIT_0 = 16'h0000;

ROM16 rom16_inst_846 (
    .DO(rom16_inst_846_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_846.INIT_0 = 16'h0000;

ROM16 rom16_inst_847 (
    .DO(rom16_inst_847_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_847.INIT_0 = 16'h0000;

ROM16 rom16_inst_848 (
    .DO(rom16_inst_848_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_848.INIT_0 = 16'h0000;

ROM16 rom16_inst_849 (
    .DO(rom16_inst_849_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_849.INIT_0 = 16'h0000;

ROM16 rom16_inst_850 (
    .DO(rom16_inst_850_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_850.INIT_0 = 16'h0000;

ROM16 rom16_inst_851 (
    .DO(rom16_inst_851_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_851.INIT_0 = 16'h0000;

ROM16 rom16_inst_852 (
    .DO(rom16_inst_852_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_852.INIT_0 = 16'h0000;

ROM16 rom16_inst_853 (
    .DO(rom16_inst_853_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_853.INIT_0 = 16'h0000;

ROM16 rom16_inst_854 (
    .DO(rom16_inst_854_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_854.INIT_0 = 16'h0000;

ROM16 rom16_inst_855 (
    .DO(rom16_inst_855_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_855.INIT_0 = 16'h0000;

ROM16 rom16_inst_856 (
    .DO(rom16_inst_856_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_856.INIT_0 = 16'h0000;

ROM16 rom16_inst_857 (
    .DO(rom16_inst_857_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_857.INIT_0 = 16'h0000;

ROM16 rom16_inst_858 (
    .DO(rom16_inst_858_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_858.INIT_0 = 16'h0000;

ROM16 rom16_inst_859 (
    .DO(rom16_inst_859_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_859.INIT_0 = 16'h0000;

ROM16 rom16_inst_860 (
    .DO(rom16_inst_860_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_860.INIT_0 = 16'h0000;

ROM16 rom16_inst_861 (
    .DO(rom16_inst_861_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_861.INIT_0 = 16'h0000;

ROM16 rom16_inst_862 (
    .DO(rom16_inst_862_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_862.INIT_0 = 16'h0000;

ROM16 rom16_inst_863 (
    .DO(rom16_inst_863_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_863.INIT_0 = 16'h0000;

ROM16 rom16_inst_864 (
    .DO(rom16_inst_864_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_864.INIT_0 = 16'h0000;

ROM16 rom16_inst_865 (
    .DO(rom16_inst_865_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_865.INIT_0 = 16'h0000;

ROM16 rom16_inst_866 (
    .DO(rom16_inst_866_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_866.INIT_0 = 16'h0000;

ROM16 rom16_inst_867 (
    .DO(rom16_inst_867_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_867.INIT_0 = 16'h0000;

ROM16 rom16_inst_868 (
    .DO(rom16_inst_868_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_868.INIT_0 = 16'h0000;

ROM16 rom16_inst_869 (
    .DO(rom16_inst_869_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_869.INIT_0 = 16'h0000;

ROM16 rom16_inst_870 (
    .DO(rom16_inst_870_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_870.INIT_0 = 16'h0000;

ROM16 rom16_inst_871 (
    .DO(rom16_inst_871_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_871.INIT_0 = 16'h0000;

ROM16 rom16_inst_872 (
    .DO(rom16_inst_872_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_872.INIT_0 = 16'h0000;

ROM16 rom16_inst_873 (
    .DO(rom16_inst_873_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_873.INIT_0 = 16'h0000;

ROM16 rom16_inst_874 (
    .DO(rom16_inst_874_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_874.INIT_0 = 16'h0000;

ROM16 rom16_inst_875 (
    .DO(rom16_inst_875_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_875.INIT_0 = 16'h0000;

ROM16 rom16_inst_876 (
    .DO(rom16_inst_876_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_876.INIT_0 = 16'h0000;

ROM16 rom16_inst_877 (
    .DO(rom16_inst_877_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_877.INIT_0 = 16'h0000;

ROM16 rom16_inst_878 (
    .DO(rom16_inst_878_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_878.INIT_0 = 16'h0000;

ROM16 rom16_inst_879 (
    .DO(rom16_inst_879_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_879.INIT_0 = 16'h0000;

ROM16 rom16_inst_880 (
    .DO(rom16_inst_880_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_880.INIT_0 = 16'h0000;

ROM16 rom16_inst_881 (
    .DO(rom16_inst_881_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_881.INIT_0 = 16'h0000;

ROM16 rom16_inst_882 (
    .DO(rom16_inst_882_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_882.INIT_0 = 16'h0000;

ROM16 rom16_inst_883 (
    .DO(rom16_inst_883_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_883.INIT_0 = 16'h0000;

ROM16 rom16_inst_884 (
    .DO(rom16_inst_884_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_884.INIT_0 = 16'h0000;

ROM16 rom16_inst_885 (
    .DO(rom16_inst_885_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_885.INIT_0 = 16'h0000;

ROM16 rom16_inst_886 (
    .DO(rom16_inst_886_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_886.INIT_0 = 16'h0000;

ROM16 rom16_inst_887 (
    .DO(rom16_inst_887_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_887.INIT_0 = 16'h0000;

ROM16 rom16_inst_888 (
    .DO(rom16_inst_888_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_888.INIT_0 = 16'h0000;

ROM16 rom16_inst_889 (
    .DO(rom16_inst_889_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_889.INIT_0 = 16'h0000;

ROM16 rom16_inst_890 (
    .DO(rom16_inst_890_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_890.INIT_0 = 16'h0000;

ROM16 rom16_inst_891 (
    .DO(rom16_inst_891_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_891.INIT_0 = 16'h0000;

ROM16 rom16_inst_892 (
    .DO(rom16_inst_892_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_892.INIT_0 = 16'h0000;

ROM16 rom16_inst_893 (
    .DO(rom16_inst_893_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_893.INIT_0 = 16'h0000;

ROM16 rom16_inst_894 (
    .DO(rom16_inst_894_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_894.INIT_0 = 16'h0000;

ROM16 rom16_inst_895 (
    .DO(rom16_inst_895_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_895.INIT_0 = 16'h0000;

ROM16 rom16_inst_896 (
    .DO(rom16_inst_896_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_896.INIT_0 = 16'h0000;

ROM16 rom16_inst_897 (
    .DO(rom16_inst_897_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_897.INIT_0 = 16'h0000;

ROM16 rom16_inst_898 (
    .DO(rom16_inst_898_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_898.INIT_0 = 16'h0000;

ROM16 rom16_inst_899 (
    .DO(rom16_inst_899_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_899.INIT_0 = 16'h0000;

ROM16 rom16_inst_900 (
    .DO(rom16_inst_900_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_900.INIT_0 = 16'h0000;

ROM16 rom16_inst_901 (
    .DO(rom16_inst_901_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_901.INIT_0 = 16'h0000;

ROM16 rom16_inst_902 (
    .DO(rom16_inst_902_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_902.INIT_0 = 16'h0000;

ROM16 rom16_inst_903 (
    .DO(rom16_inst_903_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_903.INIT_0 = 16'h0000;

ROM16 rom16_inst_904 (
    .DO(rom16_inst_904_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_904.INIT_0 = 16'h0000;

ROM16 rom16_inst_905 (
    .DO(rom16_inst_905_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_905.INIT_0 = 16'h0000;

ROM16 rom16_inst_906 (
    .DO(rom16_inst_906_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_906.INIT_0 = 16'h0000;

ROM16 rom16_inst_907 (
    .DO(rom16_inst_907_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_907.INIT_0 = 16'h0000;

ROM16 rom16_inst_908 (
    .DO(rom16_inst_908_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_908.INIT_0 = 16'h0000;

ROM16 rom16_inst_909 (
    .DO(rom16_inst_909_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_909.INIT_0 = 16'h0000;

ROM16 rom16_inst_910 (
    .DO(rom16_inst_910_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_910.INIT_0 = 16'h0000;

ROM16 rom16_inst_911 (
    .DO(rom16_inst_911_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_911.INIT_0 = 16'h0000;

ROM16 rom16_inst_912 (
    .DO(rom16_inst_912_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_912.INIT_0 = 16'h0000;

ROM16 rom16_inst_913 (
    .DO(rom16_inst_913_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_913.INIT_0 = 16'h0000;

ROM16 rom16_inst_914 (
    .DO(rom16_inst_914_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_914.INIT_0 = 16'h0000;

ROM16 rom16_inst_915 (
    .DO(rom16_inst_915_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_915.INIT_0 = 16'h0000;

ROM16 rom16_inst_916 (
    .DO(rom16_inst_916_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_916.INIT_0 = 16'h0000;

ROM16 rom16_inst_917 (
    .DO(rom16_inst_917_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_917.INIT_0 = 16'h0000;

ROM16 rom16_inst_918 (
    .DO(rom16_inst_918_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_918.INIT_0 = 16'h0000;

ROM16 rom16_inst_919 (
    .DO(rom16_inst_919_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_919.INIT_0 = 16'h0000;

ROM16 rom16_inst_920 (
    .DO(rom16_inst_920_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_920.INIT_0 = 16'h0000;

ROM16 rom16_inst_921 (
    .DO(rom16_inst_921_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_921.INIT_0 = 16'h0000;

ROM16 rom16_inst_922 (
    .DO(rom16_inst_922_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_922.INIT_0 = 16'h0000;

ROM16 rom16_inst_923 (
    .DO(rom16_inst_923_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_923.INIT_0 = 16'h0000;

ROM16 rom16_inst_924 (
    .DO(rom16_inst_924_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_924.INIT_0 = 16'h0000;

ROM16 rom16_inst_925 (
    .DO(rom16_inst_925_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_925.INIT_0 = 16'h0000;

ROM16 rom16_inst_926 (
    .DO(rom16_inst_926_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_926.INIT_0 = 16'h0000;

ROM16 rom16_inst_927 (
    .DO(rom16_inst_927_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_927.INIT_0 = 16'h0000;

ROM16 rom16_inst_928 (
    .DO(rom16_inst_928_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_928.INIT_0 = 16'h0000;

ROM16 rom16_inst_929 (
    .DO(rom16_inst_929_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_929.INIT_0 = 16'h0000;

ROM16 rom16_inst_930 (
    .DO(rom16_inst_930_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_930.INIT_0 = 16'h0000;

ROM16 rom16_inst_931 (
    .DO(rom16_inst_931_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_931.INIT_0 = 16'h0000;

ROM16 rom16_inst_932 (
    .DO(rom16_inst_932_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_932.INIT_0 = 16'h0000;

ROM16 rom16_inst_933 (
    .DO(rom16_inst_933_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_933.INIT_0 = 16'h0000;

ROM16 rom16_inst_934 (
    .DO(rom16_inst_934_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_934.INIT_0 = 16'h0000;

ROM16 rom16_inst_935 (
    .DO(rom16_inst_935_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_935.INIT_0 = 16'h0000;

ROM16 rom16_inst_936 (
    .DO(rom16_inst_936_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_936.INIT_0 = 16'h0000;

ROM16 rom16_inst_937 (
    .DO(rom16_inst_937_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_937.INIT_0 = 16'h0000;

ROM16 rom16_inst_938 (
    .DO(rom16_inst_938_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_938.INIT_0 = 16'h0000;

ROM16 rom16_inst_939 (
    .DO(rom16_inst_939_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_939.INIT_0 = 16'h0000;

ROM16 rom16_inst_940 (
    .DO(rom16_inst_940_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_940.INIT_0 = 16'h0000;

ROM16 rom16_inst_941 (
    .DO(rom16_inst_941_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_941.INIT_0 = 16'h0000;

ROM16 rom16_inst_942 (
    .DO(rom16_inst_942_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_942.INIT_0 = 16'h0000;

ROM16 rom16_inst_943 (
    .DO(rom16_inst_943_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_943.INIT_0 = 16'h0000;

ROM16 rom16_inst_944 (
    .DO(rom16_inst_944_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_944.INIT_0 = 16'h0000;

ROM16 rom16_inst_945 (
    .DO(rom16_inst_945_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_945.INIT_0 = 16'h0000;

ROM16 rom16_inst_946 (
    .DO(rom16_inst_946_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_946.INIT_0 = 16'h0000;

ROM16 rom16_inst_947 (
    .DO(rom16_inst_947_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_947.INIT_0 = 16'h0000;

ROM16 rom16_inst_948 (
    .DO(rom16_inst_948_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_948.INIT_0 = 16'h0000;

ROM16 rom16_inst_949 (
    .DO(rom16_inst_949_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_949.INIT_0 = 16'h0000;

ROM16 rom16_inst_950 (
    .DO(rom16_inst_950_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_950.INIT_0 = 16'h0000;

ROM16 rom16_inst_951 (
    .DO(rom16_inst_951_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_951.INIT_0 = 16'h0000;

ROM16 rom16_inst_952 (
    .DO(rom16_inst_952_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_952.INIT_0 = 16'h0000;

ROM16 rom16_inst_953 (
    .DO(rom16_inst_953_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_953.INIT_0 = 16'h0000;

ROM16 rom16_inst_954 (
    .DO(rom16_inst_954_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_954.INIT_0 = 16'h0000;

ROM16 rom16_inst_955 (
    .DO(rom16_inst_955_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_955.INIT_0 = 16'h0000;

ROM16 rom16_inst_956 (
    .DO(rom16_inst_956_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_956.INIT_0 = 16'h0000;

ROM16 rom16_inst_957 (
    .DO(rom16_inst_957_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_957.INIT_0 = 16'h0000;

ROM16 rom16_inst_958 (
    .DO(rom16_inst_958_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_958.INIT_0 = 16'h0000;

ROM16 rom16_inst_959 (
    .DO(rom16_inst_959_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_959.INIT_0 = 16'h0000;

ROM16 rom16_inst_960 (
    .DO(rom16_inst_960_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_960.INIT_0 = 16'h0000;

ROM16 rom16_inst_961 (
    .DO(rom16_inst_961_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_961.INIT_0 = 16'h0000;

ROM16 rom16_inst_962 (
    .DO(rom16_inst_962_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_962.INIT_0 = 16'h0000;

ROM16 rom16_inst_963 (
    .DO(rom16_inst_963_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_963.INIT_0 = 16'h0000;

ROM16 rom16_inst_964 (
    .DO(rom16_inst_964_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_964.INIT_0 = 16'h0000;

ROM16 rom16_inst_965 (
    .DO(rom16_inst_965_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_965.INIT_0 = 16'h0000;

ROM16 rom16_inst_966 (
    .DO(rom16_inst_966_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_966.INIT_0 = 16'h0000;

ROM16 rom16_inst_967 (
    .DO(rom16_inst_967_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_967.INIT_0 = 16'h0000;

ROM16 rom16_inst_968 (
    .DO(rom16_inst_968_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_968.INIT_0 = 16'h0000;

ROM16 rom16_inst_969 (
    .DO(rom16_inst_969_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_969.INIT_0 = 16'h0000;

ROM16 rom16_inst_970 (
    .DO(rom16_inst_970_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_970.INIT_0 = 16'h0000;

ROM16 rom16_inst_971 (
    .DO(rom16_inst_971_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_971.INIT_0 = 16'h0000;

ROM16 rom16_inst_972 (
    .DO(rom16_inst_972_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_972.INIT_0 = 16'h0000;

ROM16 rom16_inst_973 (
    .DO(rom16_inst_973_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_973.INIT_0 = 16'h0000;

ROM16 rom16_inst_974 (
    .DO(rom16_inst_974_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_974.INIT_0 = 16'h0000;

ROM16 rom16_inst_975 (
    .DO(rom16_inst_975_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_975.INIT_0 = 16'h0000;

ROM16 rom16_inst_976 (
    .DO(rom16_inst_976_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_976.INIT_0 = 16'h0000;

ROM16 rom16_inst_977 (
    .DO(rom16_inst_977_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_977.INIT_0 = 16'h0000;

ROM16 rom16_inst_978 (
    .DO(rom16_inst_978_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_978.INIT_0 = 16'h0000;

ROM16 rom16_inst_979 (
    .DO(rom16_inst_979_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_979.INIT_0 = 16'h0000;

ROM16 rom16_inst_980 (
    .DO(rom16_inst_980_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_980.INIT_0 = 16'h0000;

ROM16 rom16_inst_981 (
    .DO(rom16_inst_981_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_981.INIT_0 = 16'h0000;

ROM16 rom16_inst_982 (
    .DO(rom16_inst_982_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_982.INIT_0 = 16'h0000;

ROM16 rom16_inst_983 (
    .DO(rom16_inst_983_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_983.INIT_0 = 16'h0000;

ROM16 rom16_inst_984 (
    .DO(rom16_inst_984_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_984.INIT_0 = 16'h0000;

ROM16 rom16_inst_985 (
    .DO(rom16_inst_985_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_985.INIT_0 = 16'h0000;

ROM16 rom16_inst_986 (
    .DO(rom16_inst_986_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_986.INIT_0 = 16'h0000;

ROM16 rom16_inst_987 (
    .DO(rom16_inst_987_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_987.INIT_0 = 16'h0000;

ROM16 rom16_inst_988 (
    .DO(rom16_inst_988_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_988.INIT_0 = 16'h0000;

ROM16 rom16_inst_989 (
    .DO(rom16_inst_989_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_989.INIT_0 = 16'h0000;

ROM16 rom16_inst_990 (
    .DO(rom16_inst_990_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_990.INIT_0 = 16'h0000;

ROM16 rom16_inst_991 (
    .DO(rom16_inst_991_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_991.INIT_0 = 16'h0000;

ROM16 rom16_inst_992 (
    .DO(rom16_inst_992_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_992.INIT_0 = 16'h0000;

ROM16 rom16_inst_993 (
    .DO(rom16_inst_993_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_993.INIT_0 = 16'h0000;

ROM16 rom16_inst_994 (
    .DO(rom16_inst_994_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_994.INIT_0 = 16'h0000;

ROM16 rom16_inst_995 (
    .DO(rom16_inst_995_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_995.INIT_0 = 16'h0000;

ROM16 rom16_inst_996 (
    .DO(rom16_inst_996_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_996.INIT_0 = 16'h0000;

ROM16 rom16_inst_997 (
    .DO(rom16_inst_997_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_997.INIT_0 = 16'h0000;

ROM16 rom16_inst_998 (
    .DO(rom16_inst_998_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_998.INIT_0 = 16'h0000;

ROM16 rom16_inst_999 (
    .DO(rom16_inst_999_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_999.INIT_0 = 16'h0000;

ROM16 rom16_inst_1000 (
    .DO(rom16_inst_1000_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_1000.INIT_0 = 16'h0000;

ROM16 rom16_inst_1001 (
    .DO(rom16_inst_1001_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_1001.INIT_0 = 16'h0000;

ROM16 rom16_inst_1002 (
    .DO(rom16_inst_1002_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_1002.INIT_0 = 16'h0000;

ROM16 rom16_inst_1003 (
    .DO(rom16_inst_1003_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_1003.INIT_0 = 16'h0000;

ROM16 rom16_inst_1004 (
    .DO(rom16_inst_1004_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_1004.INIT_0 = 16'h0000;

ROM16 rom16_inst_1005 (
    .DO(rom16_inst_1005_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_1005.INIT_0 = 16'h0000;

ROM16 rom16_inst_1006 (
    .DO(rom16_inst_1006_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_1006.INIT_0 = 16'h0000;

ROM16 rom16_inst_1007 (
    .DO(rom16_inst_1007_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_1007.INIT_0 = 16'h0000;

ROM16 rom16_inst_1008 (
    .DO(rom16_inst_1008_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_1008.INIT_0 = 16'h0000;

ROM16 rom16_inst_1009 (
    .DO(rom16_inst_1009_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_1009.INIT_0 = 16'h0000;

ROM16 rom16_inst_1010 (
    .DO(rom16_inst_1010_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_1010.INIT_0 = 16'h0000;

ROM16 rom16_inst_1011 (
    .DO(rom16_inst_1011_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_1011.INIT_0 = 16'h0000;

ROM16 rom16_inst_1012 (
    .DO(rom16_inst_1012_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_1012.INIT_0 = 16'h0000;

ROM16 rom16_inst_1013 (
    .DO(rom16_inst_1013_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_1013.INIT_0 = 16'h0000;

ROM16 rom16_inst_1014 (
    .DO(rom16_inst_1014_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_1014.INIT_0 = 16'h0000;

ROM16 rom16_inst_1015 (
    .DO(rom16_inst_1015_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_1015.INIT_0 = 16'h0000;

ROM16 rom16_inst_1016 (
    .DO(rom16_inst_1016_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_1016.INIT_0 = 16'h0000;

ROM16 rom16_inst_1017 (
    .DO(rom16_inst_1017_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_1017.INIT_0 = 16'h0000;

ROM16 rom16_inst_1018 (
    .DO(rom16_inst_1018_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_1018.INIT_0 = 16'h0000;

ROM16 rom16_inst_1019 (
    .DO(rom16_inst_1019_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_1019.INIT_0 = 16'h0000;

ROM16 rom16_inst_1020 (
    .DO(rom16_inst_1020_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_1020.INIT_0 = 16'h0000;

ROM16 rom16_inst_1021 (
    .DO(rom16_inst_1021_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_1021.INIT_0 = 16'h0000;

ROM16 rom16_inst_1022 (
    .DO(rom16_inst_1022_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_1022.INIT_0 = 16'h0000;

ROM16 rom16_inst_1023 (
    .DO(rom16_inst_1023_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_1023.INIT_0 = 16'h0000;

MUX2 mux_inst_0 (
  .O(mux_o_0),
  .I0(rom16_inst_0_dout[0]),
  .I1(rom16_inst_16_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_1 (
  .O(mux_o_1),
  .I0(rom16_inst_32_dout[0]),
  .I1(rom16_inst_48_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_2 (
  .O(mux_o_2),
  .I0(rom16_inst_64_dout[0]),
  .I1(rom16_inst_80_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_3 (
  .O(mux_o_3),
  .I0(rom16_inst_96_dout[0]),
  .I1(rom16_inst_112_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_4 (
  .O(mux_o_4),
  .I0(rom16_inst_128_dout[0]),
  .I1(rom16_inst_144_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_5 (
  .O(mux_o_5),
  .I0(rom16_inst_160_dout[0]),
  .I1(rom16_inst_176_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_6 (
  .O(mux_o_6),
  .I0(rom16_inst_192_dout[0]),
  .I1(rom16_inst_208_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_7 (
  .O(mux_o_7),
  .I0(rom16_inst_224_dout[0]),
  .I1(rom16_inst_240_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_8 (
  .O(mux_o_8),
  .I0(rom16_inst_256_dout[0]),
  .I1(rom16_inst_272_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_9 (
  .O(mux_o_9),
  .I0(rom16_inst_288_dout[0]),
  .I1(rom16_inst_304_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_10 (
  .O(mux_o_10),
  .I0(rom16_inst_320_dout[0]),
  .I1(rom16_inst_336_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_11 (
  .O(mux_o_11),
  .I0(rom16_inst_352_dout[0]),
  .I1(rom16_inst_368_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_12 (
  .O(mux_o_12),
  .I0(rom16_inst_384_dout[0]),
  .I1(rom16_inst_400_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_13 (
  .O(mux_o_13),
  .I0(rom16_inst_416_dout[0]),
  .I1(rom16_inst_432_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_14 (
  .O(mux_o_14),
  .I0(rom16_inst_448_dout[0]),
  .I1(rom16_inst_464_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_15 (
  .O(mux_o_15),
  .I0(rom16_inst_480_dout[0]),
  .I1(rom16_inst_496_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_16 (
  .O(mux_o_16),
  .I0(rom16_inst_512_dout[0]),
  .I1(rom16_inst_528_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_17 (
  .O(mux_o_17),
  .I0(rom16_inst_544_dout[0]),
  .I1(rom16_inst_560_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_18 (
  .O(mux_o_18),
  .I0(rom16_inst_576_dout[0]),
  .I1(rom16_inst_592_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_19 (
  .O(mux_o_19),
  .I0(rom16_inst_608_dout[0]),
  .I1(rom16_inst_624_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_20 (
  .O(mux_o_20),
  .I0(rom16_inst_640_dout[0]),
  .I1(rom16_inst_656_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_21 (
  .O(mux_o_21),
  .I0(rom16_inst_672_dout[0]),
  .I1(rom16_inst_688_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_22 (
  .O(mux_o_22),
  .I0(rom16_inst_704_dout[0]),
  .I1(rom16_inst_720_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_23 (
  .O(mux_o_23),
  .I0(rom16_inst_736_dout[0]),
  .I1(rom16_inst_752_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_24 (
  .O(mux_o_24),
  .I0(rom16_inst_768_dout[0]),
  .I1(rom16_inst_784_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_25 (
  .O(mux_o_25),
  .I0(rom16_inst_800_dout[0]),
  .I1(rom16_inst_816_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_26 (
  .O(mux_o_26),
  .I0(rom16_inst_832_dout[0]),
  .I1(rom16_inst_848_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_27 (
  .O(mux_o_27),
  .I0(rom16_inst_864_dout[0]),
  .I1(rom16_inst_880_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_28 (
  .O(mux_o_28),
  .I0(rom16_inst_896_dout[0]),
  .I1(rom16_inst_912_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_29 (
  .O(mux_o_29),
  .I0(rom16_inst_928_dout[0]),
  .I1(rom16_inst_944_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_30 (
  .O(mux_o_30),
  .I0(rom16_inst_960_dout[0]),
  .I1(rom16_inst_976_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_31 (
  .O(mux_o_31),
  .I0(rom16_inst_992_dout[0]),
  .I1(rom16_inst_1008_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_32 (
  .O(mux_o_32),
  .I0(mux_o_0),
  .I1(mux_o_1),
  .S0(ad[5])
);
MUX2 mux_inst_33 (
  .O(mux_o_33),
  .I0(mux_o_2),
  .I1(mux_o_3),
  .S0(ad[5])
);
MUX2 mux_inst_34 (
  .O(mux_o_34),
  .I0(mux_o_4),
  .I1(mux_o_5),
  .S0(ad[5])
);
MUX2 mux_inst_35 (
  .O(mux_o_35),
  .I0(mux_o_6),
  .I1(mux_o_7),
  .S0(ad[5])
);
MUX2 mux_inst_36 (
  .O(mux_o_36),
  .I0(mux_o_8),
  .I1(mux_o_9),
  .S0(ad[5])
);
MUX2 mux_inst_37 (
  .O(mux_o_37),
  .I0(mux_o_10),
  .I1(mux_o_11),
  .S0(ad[5])
);
MUX2 mux_inst_38 (
  .O(mux_o_38),
  .I0(mux_o_12),
  .I1(mux_o_13),
  .S0(ad[5])
);
MUX2 mux_inst_39 (
  .O(mux_o_39),
  .I0(mux_o_14),
  .I1(mux_o_15),
  .S0(ad[5])
);
MUX2 mux_inst_40 (
  .O(mux_o_40),
  .I0(mux_o_16),
  .I1(mux_o_17),
  .S0(ad[5])
);
MUX2 mux_inst_41 (
  .O(mux_o_41),
  .I0(mux_o_18),
  .I1(mux_o_19),
  .S0(ad[5])
);
MUX2 mux_inst_42 (
  .O(mux_o_42),
  .I0(mux_o_20),
  .I1(mux_o_21),
  .S0(ad[5])
);
MUX2 mux_inst_43 (
  .O(mux_o_43),
  .I0(mux_o_22),
  .I1(mux_o_23),
  .S0(ad[5])
);
MUX2 mux_inst_44 (
  .O(mux_o_44),
  .I0(mux_o_24),
  .I1(mux_o_25),
  .S0(ad[5])
);
MUX2 mux_inst_45 (
  .O(mux_o_45),
  .I0(mux_o_26),
  .I1(mux_o_27),
  .S0(ad[5])
);
MUX2 mux_inst_46 (
  .O(mux_o_46),
  .I0(mux_o_28),
  .I1(mux_o_29),
  .S0(ad[5])
);
MUX2 mux_inst_47 (
  .O(mux_o_47),
  .I0(mux_o_30),
  .I1(mux_o_31),
  .S0(ad[5])
);
MUX2 mux_inst_48 (
  .O(mux_o_48),
  .I0(mux_o_32),
  .I1(mux_o_33),
  .S0(ad[6])
);
MUX2 mux_inst_49 (
  .O(mux_o_49),
  .I0(mux_o_34),
  .I1(mux_o_35),
  .S0(ad[6])
);
MUX2 mux_inst_50 (
  .O(mux_o_50),
  .I0(mux_o_36),
  .I1(mux_o_37),
  .S0(ad[6])
);
MUX2 mux_inst_51 (
  .O(mux_o_51),
  .I0(mux_o_38),
  .I1(mux_o_39),
  .S0(ad[6])
);
MUX2 mux_inst_52 (
  .O(mux_o_52),
  .I0(mux_o_40),
  .I1(mux_o_41),
  .S0(ad[6])
);
MUX2 mux_inst_53 (
  .O(mux_o_53),
  .I0(mux_o_42),
  .I1(mux_o_43),
  .S0(ad[6])
);
MUX2 mux_inst_54 (
  .O(mux_o_54),
  .I0(mux_o_44),
  .I1(mux_o_45),
  .S0(ad[6])
);
MUX2 mux_inst_55 (
  .O(mux_o_55),
  .I0(mux_o_46),
  .I1(mux_o_47),
  .S0(ad[6])
);
MUX2 mux_inst_56 (
  .O(mux_o_56),
  .I0(mux_o_48),
  .I1(mux_o_49),
  .S0(ad[7])
);
MUX2 mux_inst_57 (
  .O(mux_o_57),
  .I0(mux_o_50),
  .I1(mux_o_51),
  .S0(ad[7])
);
MUX2 mux_inst_58 (
  .O(mux_o_58),
  .I0(mux_o_52),
  .I1(mux_o_53),
  .S0(ad[7])
);
MUX2 mux_inst_59 (
  .O(mux_o_59),
  .I0(mux_o_54),
  .I1(mux_o_55),
  .S0(ad[7])
);
MUX2 mux_inst_60 (
  .O(mux_o_60),
  .I0(mux_o_56),
  .I1(mux_o_57),
  .S0(ad[8])
);
MUX2 mux_inst_61 (
  .O(mux_o_61),
  .I0(mux_o_58),
  .I1(mux_o_59),
  .S0(ad[8])
);
MUX2 mux_inst_62 (
  .O(dout[0]),
  .I0(mux_o_60),
  .I1(mux_o_61),
  .S0(ad[9])
);
MUX2 mux_inst_63 (
  .O(mux_o_63),
  .I0(rom16_inst_1_dout[1]),
  .I1(rom16_inst_17_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_64 (
  .O(mux_o_64),
  .I0(rom16_inst_33_dout[1]),
  .I1(rom16_inst_49_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_65 (
  .O(mux_o_65),
  .I0(rom16_inst_65_dout[1]),
  .I1(rom16_inst_81_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_66 (
  .O(mux_o_66),
  .I0(rom16_inst_97_dout[1]),
  .I1(rom16_inst_113_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_67 (
  .O(mux_o_67),
  .I0(rom16_inst_129_dout[1]),
  .I1(rom16_inst_145_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_68 (
  .O(mux_o_68),
  .I0(rom16_inst_161_dout[1]),
  .I1(rom16_inst_177_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_69 (
  .O(mux_o_69),
  .I0(rom16_inst_193_dout[1]),
  .I1(rom16_inst_209_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_70 (
  .O(mux_o_70),
  .I0(rom16_inst_225_dout[1]),
  .I1(rom16_inst_241_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_71 (
  .O(mux_o_71),
  .I0(rom16_inst_257_dout[1]),
  .I1(rom16_inst_273_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_72 (
  .O(mux_o_72),
  .I0(rom16_inst_289_dout[1]),
  .I1(rom16_inst_305_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_73 (
  .O(mux_o_73),
  .I0(rom16_inst_321_dout[1]),
  .I1(rom16_inst_337_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_74 (
  .O(mux_o_74),
  .I0(rom16_inst_353_dout[1]),
  .I1(rom16_inst_369_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_75 (
  .O(mux_o_75),
  .I0(rom16_inst_385_dout[1]),
  .I1(rom16_inst_401_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_76 (
  .O(mux_o_76),
  .I0(rom16_inst_417_dout[1]),
  .I1(rom16_inst_433_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_77 (
  .O(mux_o_77),
  .I0(rom16_inst_449_dout[1]),
  .I1(rom16_inst_465_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_78 (
  .O(mux_o_78),
  .I0(rom16_inst_481_dout[1]),
  .I1(rom16_inst_497_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_79 (
  .O(mux_o_79),
  .I0(rom16_inst_513_dout[1]),
  .I1(rom16_inst_529_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_80 (
  .O(mux_o_80),
  .I0(rom16_inst_545_dout[1]),
  .I1(rom16_inst_561_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_81 (
  .O(mux_o_81),
  .I0(rom16_inst_577_dout[1]),
  .I1(rom16_inst_593_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_82 (
  .O(mux_o_82),
  .I0(rom16_inst_609_dout[1]),
  .I1(rom16_inst_625_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_83 (
  .O(mux_o_83),
  .I0(rom16_inst_641_dout[1]),
  .I1(rom16_inst_657_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_84 (
  .O(mux_o_84),
  .I0(rom16_inst_673_dout[1]),
  .I1(rom16_inst_689_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_85 (
  .O(mux_o_85),
  .I0(rom16_inst_705_dout[1]),
  .I1(rom16_inst_721_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_86 (
  .O(mux_o_86),
  .I0(rom16_inst_737_dout[1]),
  .I1(rom16_inst_753_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_87 (
  .O(mux_o_87),
  .I0(rom16_inst_769_dout[1]),
  .I1(rom16_inst_785_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_88 (
  .O(mux_o_88),
  .I0(rom16_inst_801_dout[1]),
  .I1(rom16_inst_817_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_89 (
  .O(mux_o_89),
  .I0(rom16_inst_833_dout[1]),
  .I1(rom16_inst_849_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_90 (
  .O(mux_o_90),
  .I0(rom16_inst_865_dout[1]),
  .I1(rom16_inst_881_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_91 (
  .O(mux_o_91),
  .I0(rom16_inst_897_dout[1]),
  .I1(rom16_inst_913_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_92 (
  .O(mux_o_92),
  .I0(rom16_inst_929_dout[1]),
  .I1(rom16_inst_945_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_93 (
  .O(mux_o_93),
  .I0(rom16_inst_961_dout[1]),
  .I1(rom16_inst_977_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_94 (
  .O(mux_o_94),
  .I0(rom16_inst_993_dout[1]),
  .I1(rom16_inst_1009_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_95 (
  .O(mux_o_95),
  .I0(mux_o_63),
  .I1(mux_o_64),
  .S0(ad[5])
);
MUX2 mux_inst_96 (
  .O(mux_o_96),
  .I0(mux_o_65),
  .I1(mux_o_66),
  .S0(ad[5])
);
MUX2 mux_inst_97 (
  .O(mux_o_97),
  .I0(mux_o_67),
  .I1(mux_o_68),
  .S0(ad[5])
);
MUX2 mux_inst_98 (
  .O(mux_o_98),
  .I0(mux_o_69),
  .I1(mux_o_70),
  .S0(ad[5])
);
MUX2 mux_inst_99 (
  .O(mux_o_99),
  .I0(mux_o_71),
  .I1(mux_o_72),
  .S0(ad[5])
);
MUX2 mux_inst_100 (
  .O(mux_o_100),
  .I0(mux_o_73),
  .I1(mux_o_74),
  .S0(ad[5])
);
MUX2 mux_inst_101 (
  .O(mux_o_101),
  .I0(mux_o_75),
  .I1(mux_o_76),
  .S0(ad[5])
);
MUX2 mux_inst_102 (
  .O(mux_o_102),
  .I0(mux_o_77),
  .I1(mux_o_78),
  .S0(ad[5])
);
MUX2 mux_inst_103 (
  .O(mux_o_103),
  .I0(mux_o_79),
  .I1(mux_o_80),
  .S0(ad[5])
);
MUX2 mux_inst_104 (
  .O(mux_o_104),
  .I0(mux_o_81),
  .I1(mux_o_82),
  .S0(ad[5])
);
MUX2 mux_inst_105 (
  .O(mux_o_105),
  .I0(mux_o_83),
  .I1(mux_o_84),
  .S0(ad[5])
);
MUX2 mux_inst_106 (
  .O(mux_o_106),
  .I0(mux_o_85),
  .I1(mux_o_86),
  .S0(ad[5])
);
MUX2 mux_inst_107 (
  .O(mux_o_107),
  .I0(mux_o_87),
  .I1(mux_o_88),
  .S0(ad[5])
);
MUX2 mux_inst_108 (
  .O(mux_o_108),
  .I0(mux_o_89),
  .I1(mux_o_90),
  .S0(ad[5])
);
MUX2 mux_inst_109 (
  .O(mux_o_109),
  .I0(mux_o_91),
  .I1(mux_o_92),
  .S0(ad[5])
);
MUX2 mux_inst_110 (
  .O(mux_o_110),
  .I0(mux_o_93),
  .I1(mux_o_94),
  .S0(ad[5])
);
MUX2 mux_inst_111 (
  .O(mux_o_111),
  .I0(mux_o_95),
  .I1(mux_o_96),
  .S0(ad[6])
);
MUX2 mux_inst_112 (
  .O(mux_o_112),
  .I0(mux_o_97),
  .I1(mux_o_98),
  .S0(ad[6])
);
MUX2 mux_inst_113 (
  .O(mux_o_113),
  .I0(mux_o_99),
  .I1(mux_o_100),
  .S0(ad[6])
);
MUX2 mux_inst_114 (
  .O(mux_o_114),
  .I0(mux_o_101),
  .I1(mux_o_102),
  .S0(ad[6])
);
MUX2 mux_inst_115 (
  .O(mux_o_115),
  .I0(mux_o_103),
  .I1(mux_o_104),
  .S0(ad[6])
);
MUX2 mux_inst_116 (
  .O(mux_o_116),
  .I0(mux_o_105),
  .I1(mux_o_106),
  .S0(ad[6])
);
MUX2 mux_inst_117 (
  .O(mux_o_117),
  .I0(mux_o_107),
  .I1(mux_o_108),
  .S0(ad[6])
);
MUX2 mux_inst_118 (
  .O(mux_o_118),
  .I0(mux_o_109),
  .I1(mux_o_110),
  .S0(ad[6])
);
MUX2 mux_inst_119 (
  .O(mux_o_119),
  .I0(mux_o_111),
  .I1(mux_o_112),
  .S0(ad[7])
);
MUX2 mux_inst_120 (
  .O(mux_o_120),
  .I0(mux_o_113),
  .I1(mux_o_114),
  .S0(ad[7])
);
MUX2 mux_inst_121 (
  .O(mux_o_121),
  .I0(mux_o_115),
  .I1(mux_o_116),
  .S0(ad[7])
);
MUX2 mux_inst_122 (
  .O(mux_o_122),
  .I0(mux_o_117),
  .I1(mux_o_118),
  .S0(ad[7])
);
MUX2 mux_inst_123 (
  .O(mux_o_123),
  .I0(mux_o_119),
  .I1(mux_o_120),
  .S0(ad[8])
);
MUX2 mux_inst_124 (
  .O(mux_o_124),
  .I0(mux_o_121),
  .I1(mux_o_122),
  .S0(ad[8])
);
MUX2 mux_inst_125 (
  .O(dout[1]),
  .I0(mux_o_123),
  .I1(mux_o_124),
  .S0(ad[9])
);
MUX2 mux_inst_126 (
  .O(mux_o_126),
  .I0(rom16_inst_2_dout[2]),
  .I1(rom16_inst_18_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_127 (
  .O(mux_o_127),
  .I0(rom16_inst_34_dout[2]),
  .I1(rom16_inst_50_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_128 (
  .O(mux_o_128),
  .I0(rom16_inst_66_dout[2]),
  .I1(rom16_inst_82_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_129 (
  .O(mux_o_129),
  .I0(rom16_inst_98_dout[2]),
  .I1(rom16_inst_114_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_130 (
  .O(mux_o_130),
  .I0(rom16_inst_130_dout[2]),
  .I1(rom16_inst_146_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_131 (
  .O(mux_o_131),
  .I0(rom16_inst_162_dout[2]),
  .I1(rom16_inst_178_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_132 (
  .O(mux_o_132),
  .I0(rom16_inst_194_dout[2]),
  .I1(rom16_inst_210_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_133 (
  .O(mux_o_133),
  .I0(rom16_inst_226_dout[2]),
  .I1(rom16_inst_242_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_134 (
  .O(mux_o_134),
  .I0(rom16_inst_258_dout[2]),
  .I1(rom16_inst_274_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_135 (
  .O(mux_o_135),
  .I0(rom16_inst_290_dout[2]),
  .I1(rom16_inst_306_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_136 (
  .O(mux_o_136),
  .I0(rom16_inst_322_dout[2]),
  .I1(rom16_inst_338_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_137 (
  .O(mux_o_137),
  .I0(rom16_inst_354_dout[2]),
  .I1(rom16_inst_370_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_138 (
  .O(mux_o_138),
  .I0(rom16_inst_386_dout[2]),
  .I1(rom16_inst_402_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_139 (
  .O(mux_o_139),
  .I0(rom16_inst_418_dout[2]),
  .I1(rom16_inst_434_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_140 (
  .O(mux_o_140),
  .I0(rom16_inst_450_dout[2]),
  .I1(rom16_inst_466_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_141 (
  .O(mux_o_141),
  .I0(rom16_inst_482_dout[2]),
  .I1(rom16_inst_498_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_142 (
  .O(mux_o_142),
  .I0(rom16_inst_514_dout[2]),
  .I1(rom16_inst_530_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_143 (
  .O(mux_o_143),
  .I0(rom16_inst_546_dout[2]),
  .I1(rom16_inst_562_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_144 (
  .O(mux_o_144),
  .I0(rom16_inst_578_dout[2]),
  .I1(rom16_inst_594_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_145 (
  .O(mux_o_145),
  .I0(rom16_inst_610_dout[2]),
  .I1(rom16_inst_626_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_146 (
  .O(mux_o_146),
  .I0(rom16_inst_642_dout[2]),
  .I1(rom16_inst_658_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_147 (
  .O(mux_o_147),
  .I0(rom16_inst_674_dout[2]),
  .I1(rom16_inst_690_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_148 (
  .O(mux_o_148),
  .I0(rom16_inst_706_dout[2]),
  .I1(rom16_inst_722_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_149 (
  .O(mux_o_149),
  .I0(rom16_inst_738_dout[2]),
  .I1(rom16_inst_754_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_150 (
  .O(mux_o_150),
  .I0(rom16_inst_770_dout[2]),
  .I1(rom16_inst_786_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_151 (
  .O(mux_o_151),
  .I0(rom16_inst_802_dout[2]),
  .I1(rom16_inst_818_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_152 (
  .O(mux_o_152),
  .I0(rom16_inst_834_dout[2]),
  .I1(rom16_inst_850_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_153 (
  .O(mux_o_153),
  .I0(rom16_inst_866_dout[2]),
  .I1(rom16_inst_882_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_154 (
  .O(mux_o_154),
  .I0(rom16_inst_898_dout[2]),
  .I1(rom16_inst_914_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_155 (
  .O(mux_o_155),
  .I0(rom16_inst_930_dout[2]),
  .I1(rom16_inst_946_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_156 (
  .O(mux_o_156),
  .I0(rom16_inst_962_dout[2]),
  .I1(rom16_inst_978_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_157 (
  .O(mux_o_157),
  .I0(rom16_inst_994_dout[2]),
  .I1(rom16_inst_1010_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_158 (
  .O(mux_o_158),
  .I0(mux_o_126),
  .I1(mux_o_127),
  .S0(ad[5])
);
MUX2 mux_inst_159 (
  .O(mux_o_159),
  .I0(mux_o_128),
  .I1(mux_o_129),
  .S0(ad[5])
);
MUX2 mux_inst_160 (
  .O(mux_o_160),
  .I0(mux_o_130),
  .I1(mux_o_131),
  .S0(ad[5])
);
MUX2 mux_inst_161 (
  .O(mux_o_161),
  .I0(mux_o_132),
  .I1(mux_o_133),
  .S0(ad[5])
);
MUX2 mux_inst_162 (
  .O(mux_o_162),
  .I0(mux_o_134),
  .I1(mux_o_135),
  .S0(ad[5])
);
MUX2 mux_inst_163 (
  .O(mux_o_163),
  .I0(mux_o_136),
  .I1(mux_o_137),
  .S0(ad[5])
);
MUX2 mux_inst_164 (
  .O(mux_o_164),
  .I0(mux_o_138),
  .I1(mux_o_139),
  .S0(ad[5])
);
MUX2 mux_inst_165 (
  .O(mux_o_165),
  .I0(mux_o_140),
  .I1(mux_o_141),
  .S0(ad[5])
);
MUX2 mux_inst_166 (
  .O(mux_o_166),
  .I0(mux_o_142),
  .I1(mux_o_143),
  .S0(ad[5])
);
MUX2 mux_inst_167 (
  .O(mux_o_167),
  .I0(mux_o_144),
  .I1(mux_o_145),
  .S0(ad[5])
);
MUX2 mux_inst_168 (
  .O(mux_o_168),
  .I0(mux_o_146),
  .I1(mux_o_147),
  .S0(ad[5])
);
MUX2 mux_inst_169 (
  .O(mux_o_169),
  .I0(mux_o_148),
  .I1(mux_o_149),
  .S0(ad[5])
);
MUX2 mux_inst_170 (
  .O(mux_o_170),
  .I0(mux_o_150),
  .I1(mux_o_151),
  .S0(ad[5])
);
MUX2 mux_inst_171 (
  .O(mux_o_171),
  .I0(mux_o_152),
  .I1(mux_o_153),
  .S0(ad[5])
);
MUX2 mux_inst_172 (
  .O(mux_o_172),
  .I0(mux_o_154),
  .I1(mux_o_155),
  .S0(ad[5])
);
MUX2 mux_inst_173 (
  .O(mux_o_173),
  .I0(mux_o_156),
  .I1(mux_o_157),
  .S0(ad[5])
);
MUX2 mux_inst_174 (
  .O(mux_o_174),
  .I0(mux_o_158),
  .I1(mux_o_159),
  .S0(ad[6])
);
MUX2 mux_inst_175 (
  .O(mux_o_175),
  .I0(mux_o_160),
  .I1(mux_o_161),
  .S0(ad[6])
);
MUX2 mux_inst_176 (
  .O(mux_o_176),
  .I0(mux_o_162),
  .I1(mux_o_163),
  .S0(ad[6])
);
MUX2 mux_inst_177 (
  .O(mux_o_177),
  .I0(mux_o_164),
  .I1(mux_o_165),
  .S0(ad[6])
);
MUX2 mux_inst_178 (
  .O(mux_o_178),
  .I0(mux_o_166),
  .I1(mux_o_167),
  .S0(ad[6])
);
MUX2 mux_inst_179 (
  .O(mux_o_179),
  .I0(mux_o_168),
  .I1(mux_o_169),
  .S0(ad[6])
);
MUX2 mux_inst_180 (
  .O(mux_o_180),
  .I0(mux_o_170),
  .I1(mux_o_171),
  .S0(ad[6])
);
MUX2 mux_inst_181 (
  .O(mux_o_181),
  .I0(mux_o_172),
  .I1(mux_o_173),
  .S0(ad[6])
);
MUX2 mux_inst_182 (
  .O(mux_o_182),
  .I0(mux_o_174),
  .I1(mux_o_175),
  .S0(ad[7])
);
MUX2 mux_inst_183 (
  .O(mux_o_183),
  .I0(mux_o_176),
  .I1(mux_o_177),
  .S0(ad[7])
);
MUX2 mux_inst_184 (
  .O(mux_o_184),
  .I0(mux_o_178),
  .I1(mux_o_179),
  .S0(ad[7])
);
MUX2 mux_inst_185 (
  .O(mux_o_185),
  .I0(mux_o_180),
  .I1(mux_o_181),
  .S0(ad[7])
);
MUX2 mux_inst_186 (
  .O(mux_o_186),
  .I0(mux_o_182),
  .I1(mux_o_183),
  .S0(ad[8])
);
MUX2 mux_inst_187 (
  .O(mux_o_187),
  .I0(mux_o_184),
  .I1(mux_o_185),
  .S0(ad[8])
);
MUX2 mux_inst_188 (
  .O(dout[2]),
  .I0(mux_o_186),
  .I1(mux_o_187),
  .S0(ad[9])
);
MUX2 mux_inst_189 (
  .O(mux_o_189),
  .I0(rom16_inst_3_dout[3]),
  .I1(rom16_inst_19_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_190 (
  .O(mux_o_190),
  .I0(rom16_inst_35_dout[3]),
  .I1(rom16_inst_51_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_191 (
  .O(mux_o_191),
  .I0(rom16_inst_67_dout[3]),
  .I1(rom16_inst_83_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_192 (
  .O(mux_o_192),
  .I0(rom16_inst_99_dout[3]),
  .I1(rom16_inst_115_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_193 (
  .O(mux_o_193),
  .I0(rom16_inst_131_dout[3]),
  .I1(rom16_inst_147_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_194 (
  .O(mux_o_194),
  .I0(rom16_inst_163_dout[3]),
  .I1(rom16_inst_179_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_195 (
  .O(mux_o_195),
  .I0(rom16_inst_195_dout[3]),
  .I1(rom16_inst_211_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_196 (
  .O(mux_o_196),
  .I0(rom16_inst_227_dout[3]),
  .I1(rom16_inst_243_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_197 (
  .O(mux_o_197),
  .I0(rom16_inst_259_dout[3]),
  .I1(rom16_inst_275_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_198 (
  .O(mux_o_198),
  .I0(rom16_inst_291_dout[3]),
  .I1(rom16_inst_307_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_199 (
  .O(mux_o_199),
  .I0(rom16_inst_323_dout[3]),
  .I1(rom16_inst_339_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_200 (
  .O(mux_o_200),
  .I0(rom16_inst_355_dout[3]),
  .I1(rom16_inst_371_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_201 (
  .O(mux_o_201),
  .I0(rom16_inst_387_dout[3]),
  .I1(rom16_inst_403_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_202 (
  .O(mux_o_202),
  .I0(rom16_inst_419_dout[3]),
  .I1(rom16_inst_435_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_203 (
  .O(mux_o_203),
  .I0(rom16_inst_451_dout[3]),
  .I1(rom16_inst_467_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_204 (
  .O(mux_o_204),
  .I0(rom16_inst_483_dout[3]),
  .I1(rom16_inst_499_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_205 (
  .O(mux_o_205),
  .I0(rom16_inst_515_dout[3]),
  .I1(rom16_inst_531_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_206 (
  .O(mux_o_206),
  .I0(rom16_inst_547_dout[3]),
  .I1(rom16_inst_563_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_207 (
  .O(mux_o_207),
  .I0(rom16_inst_579_dout[3]),
  .I1(rom16_inst_595_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_208 (
  .O(mux_o_208),
  .I0(rom16_inst_611_dout[3]),
  .I1(rom16_inst_627_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_209 (
  .O(mux_o_209),
  .I0(rom16_inst_643_dout[3]),
  .I1(rom16_inst_659_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_210 (
  .O(mux_o_210),
  .I0(rom16_inst_675_dout[3]),
  .I1(rom16_inst_691_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_211 (
  .O(mux_o_211),
  .I0(rom16_inst_707_dout[3]),
  .I1(rom16_inst_723_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_212 (
  .O(mux_o_212),
  .I0(rom16_inst_739_dout[3]),
  .I1(rom16_inst_755_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_213 (
  .O(mux_o_213),
  .I0(rom16_inst_771_dout[3]),
  .I1(rom16_inst_787_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_214 (
  .O(mux_o_214),
  .I0(rom16_inst_803_dout[3]),
  .I1(rom16_inst_819_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_215 (
  .O(mux_o_215),
  .I0(rom16_inst_835_dout[3]),
  .I1(rom16_inst_851_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_216 (
  .O(mux_o_216),
  .I0(rom16_inst_867_dout[3]),
  .I1(rom16_inst_883_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_217 (
  .O(mux_o_217),
  .I0(rom16_inst_899_dout[3]),
  .I1(rom16_inst_915_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_218 (
  .O(mux_o_218),
  .I0(rom16_inst_931_dout[3]),
  .I1(rom16_inst_947_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_219 (
  .O(mux_o_219),
  .I0(rom16_inst_963_dout[3]),
  .I1(rom16_inst_979_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_220 (
  .O(mux_o_220),
  .I0(rom16_inst_995_dout[3]),
  .I1(rom16_inst_1011_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_221 (
  .O(mux_o_221),
  .I0(mux_o_189),
  .I1(mux_o_190),
  .S0(ad[5])
);
MUX2 mux_inst_222 (
  .O(mux_o_222),
  .I0(mux_o_191),
  .I1(mux_o_192),
  .S0(ad[5])
);
MUX2 mux_inst_223 (
  .O(mux_o_223),
  .I0(mux_o_193),
  .I1(mux_o_194),
  .S0(ad[5])
);
MUX2 mux_inst_224 (
  .O(mux_o_224),
  .I0(mux_o_195),
  .I1(mux_o_196),
  .S0(ad[5])
);
MUX2 mux_inst_225 (
  .O(mux_o_225),
  .I0(mux_o_197),
  .I1(mux_o_198),
  .S0(ad[5])
);
MUX2 mux_inst_226 (
  .O(mux_o_226),
  .I0(mux_o_199),
  .I1(mux_o_200),
  .S0(ad[5])
);
MUX2 mux_inst_227 (
  .O(mux_o_227),
  .I0(mux_o_201),
  .I1(mux_o_202),
  .S0(ad[5])
);
MUX2 mux_inst_228 (
  .O(mux_o_228),
  .I0(mux_o_203),
  .I1(mux_o_204),
  .S0(ad[5])
);
MUX2 mux_inst_229 (
  .O(mux_o_229),
  .I0(mux_o_205),
  .I1(mux_o_206),
  .S0(ad[5])
);
MUX2 mux_inst_230 (
  .O(mux_o_230),
  .I0(mux_o_207),
  .I1(mux_o_208),
  .S0(ad[5])
);
MUX2 mux_inst_231 (
  .O(mux_o_231),
  .I0(mux_o_209),
  .I1(mux_o_210),
  .S0(ad[5])
);
MUX2 mux_inst_232 (
  .O(mux_o_232),
  .I0(mux_o_211),
  .I1(mux_o_212),
  .S0(ad[5])
);
MUX2 mux_inst_233 (
  .O(mux_o_233),
  .I0(mux_o_213),
  .I1(mux_o_214),
  .S0(ad[5])
);
MUX2 mux_inst_234 (
  .O(mux_o_234),
  .I0(mux_o_215),
  .I1(mux_o_216),
  .S0(ad[5])
);
MUX2 mux_inst_235 (
  .O(mux_o_235),
  .I0(mux_o_217),
  .I1(mux_o_218),
  .S0(ad[5])
);
MUX2 mux_inst_236 (
  .O(mux_o_236),
  .I0(mux_o_219),
  .I1(mux_o_220),
  .S0(ad[5])
);
MUX2 mux_inst_237 (
  .O(mux_o_237),
  .I0(mux_o_221),
  .I1(mux_o_222),
  .S0(ad[6])
);
MUX2 mux_inst_238 (
  .O(mux_o_238),
  .I0(mux_o_223),
  .I1(mux_o_224),
  .S0(ad[6])
);
MUX2 mux_inst_239 (
  .O(mux_o_239),
  .I0(mux_o_225),
  .I1(mux_o_226),
  .S0(ad[6])
);
MUX2 mux_inst_240 (
  .O(mux_o_240),
  .I0(mux_o_227),
  .I1(mux_o_228),
  .S0(ad[6])
);
MUX2 mux_inst_241 (
  .O(mux_o_241),
  .I0(mux_o_229),
  .I1(mux_o_230),
  .S0(ad[6])
);
MUX2 mux_inst_242 (
  .O(mux_o_242),
  .I0(mux_o_231),
  .I1(mux_o_232),
  .S0(ad[6])
);
MUX2 mux_inst_243 (
  .O(mux_o_243),
  .I0(mux_o_233),
  .I1(mux_o_234),
  .S0(ad[6])
);
MUX2 mux_inst_244 (
  .O(mux_o_244),
  .I0(mux_o_235),
  .I1(mux_o_236),
  .S0(ad[6])
);
MUX2 mux_inst_245 (
  .O(mux_o_245),
  .I0(mux_o_237),
  .I1(mux_o_238),
  .S0(ad[7])
);
MUX2 mux_inst_246 (
  .O(mux_o_246),
  .I0(mux_o_239),
  .I1(mux_o_240),
  .S0(ad[7])
);
MUX2 mux_inst_247 (
  .O(mux_o_247),
  .I0(mux_o_241),
  .I1(mux_o_242),
  .S0(ad[7])
);
MUX2 mux_inst_248 (
  .O(mux_o_248),
  .I0(mux_o_243),
  .I1(mux_o_244),
  .S0(ad[7])
);
MUX2 mux_inst_249 (
  .O(mux_o_249),
  .I0(mux_o_245),
  .I1(mux_o_246),
  .S0(ad[8])
);
MUX2 mux_inst_250 (
  .O(mux_o_250),
  .I0(mux_o_247),
  .I1(mux_o_248),
  .S0(ad[8])
);
MUX2 mux_inst_251 (
  .O(dout[3]),
  .I0(mux_o_249),
  .I1(mux_o_250),
  .S0(ad[9])
);
MUX2 mux_inst_252 (
  .O(mux_o_252),
  .I0(rom16_inst_4_dout[4]),
  .I1(rom16_inst_20_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_253 (
  .O(mux_o_253),
  .I0(rom16_inst_36_dout[4]),
  .I1(rom16_inst_52_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_254 (
  .O(mux_o_254),
  .I0(rom16_inst_68_dout[4]),
  .I1(rom16_inst_84_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_255 (
  .O(mux_o_255),
  .I0(rom16_inst_100_dout[4]),
  .I1(rom16_inst_116_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_256 (
  .O(mux_o_256),
  .I0(rom16_inst_132_dout[4]),
  .I1(rom16_inst_148_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_257 (
  .O(mux_o_257),
  .I0(rom16_inst_164_dout[4]),
  .I1(rom16_inst_180_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_258 (
  .O(mux_o_258),
  .I0(rom16_inst_196_dout[4]),
  .I1(rom16_inst_212_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_259 (
  .O(mux_o_259),
  .I0(rom16_inst_228_dout[4]),
  .I1(rom16_inst_244_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_260 (
  .O(mux_o_260),
  .I0(rom16_inst_260_dout[4]),
  .I1(rom16_inst_276_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_261 (
  .O(mux_o_261),
  .I0(rom16_inst_292_dout[4]),
  .I1(rom16_inst_308_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_262 (
  .O(mux_o_262),
  .I0(rom16_inst_324_dout[4]),
  .I1(rom16_inst_340_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_263 (
  .O(mux_o_263),
  .I0(rom16_inst_356_dout[4]),
  .I1(rom16_inst_372_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_264 (
  .O(mux_o_264),
  .I0(rom16_inst_388_dout[4]),
  .I1(rom16_inst_404_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_265 (
  .O(mux_o_265),
  .I0(rom16_inst_420_dout[4]),
  .I1(rom16_inst_436_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_266 (
  .O(mux_o_266),
  .I0(rom16_inst_452_dout[4]),
  .I1(rom16_inst_468_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_267 (
  .O(mux_o_267),
  .I0(rom16_inst_484_dout[4]),
  .I1(rom16_inst_500_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_268 (
  .O(mux_o_268),
  .I0(rom16_inst_516_dout[4]),
  .I1(rom16_inst_532_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_269 (
  .O(mux_o_269),
  .I0(rom16_inst_548_dout[4]),
  .I1(rom16_inst_564_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_270 (
  .O(mux_o_270),
  .I0(rom16_inst_580_dout[4]),
  .I1(rom16_inst_596_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_271 (
  .O(mux_o_271),
  .I0(rom16_inst_612_dout[4]),
  .I1(rom16_inst_628_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_272 (
  .O(mux_o_272),
  .I0(rom16_inst_644_dout[4]),
  .I1(rom16_inst_660_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_273 (
  .O(mux_o_273),
  .I0(rom16_inst_676_dout[4]),
  .I1(rom16_inst_692_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_274 (
  .O(mux_o_274),
  .I0(rom16_inst_708_dout[4]),
  .I1(rom16_inst_724_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_275 (
  .O(mux_o_275),
  .I0(rom16_inst_740_dout[4]),
  .I1(rom16_inst_756_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_276 (
  .O(mux_o_276),
  .I0(rom16_inst_772_dout[4]),
  .I1(rom16_inst_788_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_277 (
  .O(mux_o_277),
  .I0(rom16_inst_804_dout[4]),
  .I1(rom16_inst_820_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_278 (
  .O(mux_o_278),
  .I0(rom16_inst_836_dout[4]),
  .I1(rom16_inst_852_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_279 (
  .O(mux_o_279),
  .I0(rom16_inst_868_dout[4]),
  .I1(rom16_inst_884_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_280 (
  .O(mux_o_280),
  .I0(rom16_inst_900_dout[4]),
  .I1(rom16_inst_916_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_281 (
  .O(mux_o_281),
  .I0(rom16_inst_932_dout[4]),
  .I1(rom16_inst_948_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_282 (
  .O(mux_o_282),
  .I0(rom16_inst_964_dout[4]),
  .I1(rom16_inst_980_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_283 (
  .O(mux_o_283),
  .I0(rom16_inst_996_dout[4]),
  .I1(rom16_inst_1012_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_284 (
  .O(mux_o_284),
  .I0(mux_o_252),
  .I1(mux_o_253),
  .S0(ad[5])
);
MUX2 mux_inst_285 (
  .O(mux_o_285),
  .I0(mux_o_254),
  .I1(mux_o_255),
  .S0(ad[5])
);
MUX2 mux_inst_286 (
  .O(mux_o_286),
  .I0(mux_o_256),
  .I1(mux_o_257),
  .S0(ad[5])
);
MUX2 mux_inst_287 (
  .O(mux_o_287),
  .I0(mux_o_258),
  .I1(mux_o_259),
  .S0(ad[5])
);
MUX2 mux_inst_288 (
  .O(mux_o_288),
  .I0(mux_o_260),
  .I1(mux_o_261),
  .S0(ad[5])
);
MUX2 mux_inst_289 (
  .O(mux_o_289),
  .I0(mux_o_262),
  .I1(mux_o_263),
  .S0(ad[5])
);
MUX2 mux_inst_290 (
  .O(mux_o_290),
  .I0(mux_o_264),
  .I1(mux_o_265),
  .S0(ad[5])
);
MUX2 mux_inst_291 (
  .O(mux_o_291),
  .I0(mux_o_266),
  .I1(mux_o_267),
  .S0(ad[5])
);
MUX2 mux_inst_292 (
  .O(mux_o_292),
  .I0(mux_o_268),
  .I1(mux_o_269),
  .S0(ad[5])
);
MUX2 mux_inst_293 (
  .O(mux_o_293),
  .I0(mux_o_270),
  .I1(mux_o_271),
  .S0(ad[5])
);
MUX2 mux_inst_294 (
  .O(mux_o_294),
  .I0(mux_o_272),
  .I1(mux_o_273),
  .S0(ad[5])
);
MUX2 mux_inst_295 (
  .O(mux_o_295),
  .I0(mux_o_274),
  .I1(mux_o_275),
  .S0(ad[5])
);
MUX2 mux_inst_296 (
  .O(mux_o_296),
  .I0(mux_o_276),
  .I1(mux_o_277),
  .S0(ad[5])
);
MUX2 mux_inst_297 (
  .O(mux_o_297),
  .I0(mux_o_278),
  .I1(mux_o_279),
  .S0(ad[5])
);
MUX2 mux_inst_298 (
  .O(mux_o_298),
  .I0(mux_o_280),
  .I1(mux_o_281),
  .S0(ad[5])
);
MUX2 mux_inst_299 (
  .O(mux_o_299),
  .I0(mux_o_282),
  .I1(mux_o_283),
  .S0(ad[5])
);
MUX2 mux_inst_300 (
  .O(mux_o_300),
  .I0(mux_o_284),
  .I1(mux_o_285),
  .S0(ad[6])
);
MUX2 mux_inst_301 (
  .O(mux_o_301),
  .I0(mux_o_286),
  .I1(mux_o_287),
  .S0(ad[6])
);
MUX2 mux_inst_302 (
  .O(mux_o_302),
  .I0(mux_o_288),
  .I1(mux_o_289),
  .S0(ad[6])
);
MUX2 mux_inst_303 (
  .O(mux_o_303),
  .I0(mux_o_290),
  .I1(mux_o_291),
  .S0(ad[6])
);
MUX2 mux_inst_304 (
  .O(mux_o_304),
  .I0(mux_o_292),
  .I1(mux_o_293),
  .S0(ad[6])
);
MUX2 mux_inst_305 (
  .O(mux_o_305),
  .I0(mux_o_294),
  .I1(mux_o_295),
  .S0(ad[6])
);
MUX2 mux_inst_306 (
  .O(mux_o_306),
  .I0(mux_o_296),
  .I1(mux_o_297),
  .S0(ad[6])
);
MUX2 mux_inst_307 (
  .O(mux_o_307),
  .I0(mux_o_298),
  .I1(mux_o_299),
  .S0(ad[6])
);
MUX2 mux_inst_308 (
  .O(mux_o_308),
  .I0(mux_o_300),
  .I1(mux_o_301),
  .S0(ad[7])
);
MUX2 mux_inst_309 (
  .O(mux_o_309),
  .I0(mux_o_302),
  .I1(mux_o_303),
  .S0(ad[7])
);
MUX2 mux_inst_310 (
  .O(mux_o_310),
  .I0(mux_o_304),
  .I1(mux_o_305),
  .S0(ad[7])
);
MUX2 mux_inst_311 (
  .O(mux_o_311),
  .I0(mux_o_306),
  .I1(mux_o_307),
  .S0(ad[7])
);
MUX2 mux_inst_312 (
  .O(mux_o_312),
  .I0(mux_o_308),
  .I1(mux_o_309),
  .S0(ad[8])
);
MUX2 mux_inst_313 (
  .O(mux_o_313),
  .I0(mux_o_310),
  .I1(mux_o_311),
  .S0(ad[8])
);
MUX2 mux_inst_314 (
  .O(dout[4]),
  .I0(mux_o_312),
  .I1(mux_o_313),
  .S0(ad[9])
);
MUX2 mux_inst_315 (
  .O(mux_o_315),
  .I0(rom16_inst_5_dout[5]),
  .I1(rom16_inst_21_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_316 (
  .O(mux_o_316),
  .I0(rom16_inst_37_dout[5]),
  .I1(rom16_inst_53_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_317 (
  .O(mux_o_317),
  .I0(rom16_inst_69_dout[5]),
  .I1(rom16_inst_85_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_318 (
  .O(mux_o_318),
  .I0(rom16_inst_101_dout[5]),
  .I1(rom16_inst_117_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_319 (
  .O(mux_o_319),
  .I0(rom16_inst_133_dout[5]),
  .I1(rom16_inst_149_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_320 (
  .O(mux_o_320),
  .I0(rom16_inst_165_dout[5]),
  .I1(rom16_inst_181_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_321 (
  .O(mux_o_321),
  .I0(rom16_inst_197_dout[5]),
  .I1(rom16_inst_213_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_322 (
  .O(mux_o_322),
  .I0(rom16_inst_229_dout[5]),
  .I1(rom16_inst_245_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_323 (
  .O(mux_o_323),
  .I0(rom16_inst_261_dout[5]),
  .I1(rom16_inst_277_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_324 (
  .O(mux_o_324),
  .I0(rom16_inst_293_dout[5]),
  .I1(rom16_inst_309_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_325 (
  .O(mux_o_325),
  .I0(rom16_inst_325_dout[5]),
  .I1(rom16_inst_341_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_326 (
  .O(mux_o_326),
  .I0(rom16_inst_357_dout[5]),
  .I1(rom16_inst_373_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_327 (
  .O(mux_o_327),
  .I0(rom16_inst_389_dout[5]),
  .I1(rom16_inst_405_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_328 (
  .O(mux_o_328),
  .I0(rom16_inst_421_dout[5]),
  .I1(rom16_inst_437_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_329 (
  .O(mux_o_329),
  .I0(rom16_inst_453_dout[5]),
  .I1(rom16_inst_469_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_330 (
  .O(mux_o_330),
  .I0(rom16_inst_485_dout[5]),
  .I1(rom16_inst_501_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_331 (
  .O(mux_o_331),
  .I0(rom16_inst_517_dout[5]),
  .I1(rom16_inst_533_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_332 (
  .O(mux_o_332),
  .I0(rom16_inst_549_dout[5]),
  .I1(rom16_inst_565_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_333 (
  .O(mux_o_333),
  .I0(rom16_inst_581_dout[5]),
  .I1(rom16_inst_597_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_334 (
  .O(mux_o_334),
  .I0(rom16_inst_613_dout[5]),
  .I1(rom16_inst_629_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_335 (
  .O(mux_o_335),
  .I0(rom16_inst_645_dout[5]),
  .I1(rom16_inst_661_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_336 (
  .O(mux_o_336),
  .I0(rom16_inst_677_dout[5]),
  .I1(rom16_inst_693_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_337 (
  .O(mux_o_337),
  .I0(rom16_inst_709_dout[5]),
  .I1(rom16_inst_725_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_338 (
  .O(mux_o_338),
  .I0(rom16_inst_741_dout[5]),
  .I1(rom16_inst_757_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_339 (
  .O(mux_o_339),
  .I0(rom16_inst_773_dout[5]),
  .I1(rom16_inst_789_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_340 (
  .O(mux_o_340),
  .I0(rom16_inst_805_dout[5]),
  .I1(rom16_inst_821_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_341 (
  .O(mux_o_341),
  .I0(rom16_inst_837_dout[5]),
  .I1(rom16_inst_853_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_342 (
  .O(mux_o_342),
  .I0(rom16_inst_869_dout[5]),
  .I1(rom16_inst_885_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_343 (
  .O(mux_o_343),
  .I0(rom16_inst_901_dout[5]),
  .I1(rom16_inst_917_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_344 (
  .O(mux_o_344),
  .I0(rom16_inst_933_dout[5]),
  .I1(rom16_inst_949_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_345 (
  .O(mux_o_345),
  .I0(rom16_inst_965_dout[5]),
  .I1(rom16_inst_981_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_346 (
  .O(mux_o_346),
  .I0(rom16_inst_997_dout[5]),
  .I1(rom16_inst_1013_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_347 (
  .O(mux_o_347),
  .I0(mux_o_315),
  .I1(mux_o_316),
  .S0(ad[5])
);
MUX2 mux_inst_348 (
  .O(mux_o_348),
  .I0(mux_o_317),
  .I1(mux_o_318),
  .S0(ad[5])
);
MUX2 mux_inst_349 (
  .O(mux_o_349),
  .I0(mux_o_319),
  .I1(mux_o_320),
  .S0(ad[5])
);
MUX2 mux_inst_350 (
  .O(mux_o_350),
  .I0(mux_o_321),
  .I1(mux_o_322),
  .S0(ad[5])
);
MUX2 mux_inst_351 (
  .O(mux_o_351),
  .I0(mux_o_323),
  .I1(mux_o_324),
  .S0(ad[5])
);
MUX2 mux_inst_352 (
  .O(mux_o_352),
  .I0(mux_o_325),
  .I1(mux_o_326),
  .S0(ad[5])
);
MUX2 mux_inst_353 (
  .O(mux_o_353),
  .I0(mux_o_327),
  .I1(mux_o_328),
  .S0(ad[5])
);
MUX2 mux_inst_354 (
  .O(mux_o_354),
  .I0(mux_o_329),
  .I1(mux_o_330),
  .S0(ad[5])
);
MUX2 mux_inst_355 (
  .O(mux_o_355),
  .I0(mux_o_331),
  .I1(mux_o_332),
  .S0(ad[5])
);
MUX2 mux_inst_356 (
  .O(mux_o_356),
  .I0(mux_o_333),
  .I1(mux_o_334),
  .S0(ad[5])
);
MUX2 mux_inst_357 (
  .O(mux_o_357),
  .I0(mux_o_335),
  .I1(mux_o_336),
  .S0(ad[5])
);
MUX2 mux_inst_358 (
  .O(mux_o_358),
  .I0(mux_o_337),
  .I1(mux_o_338),
  .S0(ad[5])
);
MUX2 mux_inst_359 (
  .O(mux_o_359),
  .I0(mux_o_339),
  .I1(mux_o_340),
  .S0(ad[5])
);
MUX2 mux_inst_360 (
  .O(mux_o_360),
  .I0(mux_o_341),
  .I1(mux_o_342),
  .S0(ad[5])
);
MUX2 mux_inst_361 (
  .O(mux_o_361),
  .I0(mux_o_343),
  .I1(mux_o_344),
  .S0(ad[5])
);
MUX2 mux_inst_362 (
  .O(mux_o_362),
  .I0(mux_o_345),
  .I1(mux_o_346),
  .S0(ad[5])
);
MUX2 mux_inst_363 (
  .O(mux_o_363),
  .I0(mux_o_347),
  .I1(mux_o_348),
  .S0(ad[6])
);
MUX2 mux_inst_364 (
  .O(mux_o_364),
  .I0(mux_o_349),
  .I1(mux_o_350),
  .S0(ad[6])
);
MUX2 mux_inst_365 (
  .O(mux_o_365),
  .I0(mux_o_351),
  .I1(mux_o_352),
  .S0(ad[6])
);
MUX2 mux_inst_366 (
  .O(mux_o_366),
  .I0(mux_o_353),
  .I1(mux_o_354),
  .S0(ad[6])
);
MUX2 mux_inst_367 (
  .O(mux_o_367),
  .I0(mux_o_355),
  .I1(mux_o_356),
  .S0(ad[6])
);
MUX2 mux_inst_368 (
  .O(mux_o_368),
  .I0(mux_o_357),
  .I1(mux_o_358),
  .S0(ad[6])
);
MUX2 mux_inst_369 (
  .O(mux_o_369),
  .I0(mux_o_359),
  .I1(mux_o_360),
  .S0(ad[6])
);
MUX2 mux_inst_370 (
  .O(mux_o_370),
  .I0(mux_o_361),
  .I1(mux_o_362),
  .S0(ad[6])
);
MUX2 mux_inst_371 (
  .O(mux_o_371),
  .I0(mux_o_363),
  .I1(mux_o_364),
  .S0(ad[7])
);
MUX2 mux_inst_372 (
  .O(mux_o_372),
  .I0(mux_o_365),
  .I1(mux_o_366),
  .S0(ad[7])
);
MUX2 mux_inst_373 (
  .O(mux_o_373),
  .I0(mux_o_367),
  .I1(mux_o_368),
  .S0(ad[7])
);
MUX2 mux_inst_374 (
  .O(mux_o_374),
  .I0(mux_o_369),
  .I1(mux_o_370),
  .S0(ad[7])
);
MUX2 mux_inst_375 (
  .O(mux_o_375),
  .I0(mux_o_371),
  .I1(mux_o_372),
  .S0(ad[8])
);
MUX2 mux_inst_376 (
  .O(mux_o_376),
  .I0(mux_o_373),
  .I1(mux_o_374),
  .S0(ad[8])
);
MUX2 mux_inst_377 (
  .O(dout[5]),
  .I0(mux_o_375),
  .I1(mux_o_376),
  .S0(ad[9])
);
MUX2 mux_inst_378 (
  .O(mux_o_378),
  .I0(rom16_inst_6_dout[6]),
  .I1(rom16_inst_22_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_379 (
  .O(mux_o_379),
  .I0(rom16_inst_38_dout[6]),
  .I1(rom16_inst_54_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_380 (
  .O(mux_o_380),
  .I0(rom16_inst_70_dout[6]),
  .I1(rom16_inst_86_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_381 (
  .O(mux_o_381),
  .I0(rom16_inst_102_dout[6]),
  .I1(rom16_inst_118_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_382 (
  .O(mux_o_382),
  .I0(rom16_inst_134_dout[6]),
  .I1(rom16_inst_150_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_383 (
  .O(mux_o_383),
  .I0(rom16_inst_166_dout[6]),
  .I1(rom16_inst_182_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_384 (
  .O(mux_o_384),
  .I0(rom16_inst_198_dout[6]),
  .I1(rom16_inst_214_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_385 (
  .O(mux_o_385),
  .I0(rom16_inst_230_dout[6]),
  .I1(rom16_inst_246_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_386 (
  .O(mux_o_386),
  .I0(rom16_inst_262_dout[6]),
  .I1(rom16_inst_278_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_387 (
  .O(mux_o_387),
  .I0(rom16_inst_294_dout[6]),
  .I1(rom16_inst_310_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_388 (
  .O(mux_o_388),
  .I0(rom16_inst_326_dout[6]),
  .I1(rom16_inst_342_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_389 (
  .O(mux_o_389),
  .I0(rom16_inst_358_dout[6]),
  .I1(rom16_inst_374_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_390 (
  .O(mux_o_390),
  .I0(rom16_inst_390_dout[6]),
  .I1(rom16_inst_406_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_391 (
  .O(mux_o_391),
  .I0(rom16_inst_422_dout[6]),
  .I1(rom16_inst_438_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_392 (
  .O(mux_o_392),
  .I0(rom16_inst_454_dout[6]),
  .I1(rom16_inst_470_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_393 (
  .O(mux_o_393),
  .I0(rom16_inst_486_dout[6]),
  .I1(rom16_inst_502_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_394 (
  .O(mux_o_394),
  .I0(rom16_inst_518_dout[6]),
  .I1(rom16_inst_534_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_395 (
  .O(mux_o_395),
  .I0(rom16_inst_550_dout[6]),
  .I1(rom16_inst_566_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_396 (
  .O(mux_o_396),
  .I0(rom16_inst_582_dout[6]),
  .I1(rom16_inst_598_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_397 (
  .O(mux_o_397),
  .I0(rom16_inst_614_dout[6]),
  .I1(rom16_inst_630_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_398 (
  .O(mux_o_398),
  .I0(rom16_inst_646_dout[6]),
  .I1(rom16_inst_662_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_399 (
  .O(mux_o_399),
  .I0(rom16_inst_678_dout[6]),
  .I1(rom16_inst_694_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_400 (
  .O(mux_o_400),
  .I0(rom16_inst_710_dout[6]),
  .I1(rom16_inst_726_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_401 (
  .O(mux_o_401),
  .I0(rom16_inst_742_dout[6]),
  .I1(rom16_inst_758_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_402 (
  .O(mux_o_402),
  .I0(rom16_inst_774_dout[6]),
  .I1(rom16_inst_790_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_403 (
  .O(mux_o_403),
  .I0(rom16_inst_806_dout[6]),
  .I1(rom16_inst_822_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_404 (
  .O(mux_o_404),
  .I0(rom16_inst_838_dout[6]),
  .I1(rom16_inst_854_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_405 (
  .O(mux_o_405),
  .I0(rom16_inst_870_dout[6]),
  .I1(rom16_inst_886_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_406 (
  .O(mux_o_406),
  .I0(rom16_inst_902_dout[6]),
  .I1(rom16_inst_918_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_407 (
  .O(mux_o_407),
  .I0(rom16_inst_934_dout[6]),
  .I1(rom16_inst_950_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_408 (
  .O(mux_o_408),
  .I0(rom16_inst_966_dout[6]),
  .I1(rom16_inst_982_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_409 (
  .O(mux_o_409),
  .I0(rom16_inst_998_dout[6]),
  .I1(rom16_inst_1014_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_410 (
  .O(mux_o_410),
  .I0(mux_o_378),
  .I1(mux_o_379),
  .S0(ad[5])
);
MUX2 mux_inst_411 (
  .O(mux_o_411),
  .I0(mux_o_380),
  .I1(mux_o_381),
  .S0(ad[5])
);
MUX2 mux_inst_412 (
  .O(mux_o_412),
  .I0(mux_o_382),
  .I1(mux_o_383),
  .S0(ad[5])
);
MUX2 mux_inst_413 (
  .O(mux_o_413),
  .I0(mux_o_384),
  .I1(mux_o_385),
  .S0(ad[5])
);
MUX2 mux_inst_414 (
  .O(mux_o_414),
  .I0(mux_o_386),
  .I1(mux_o_387),
  .S0(ad[5])
);
MUX2 mux_inst_415 (
  .O(mux_o_415),
  .I0(mux_o_388),
  .I1(mux_o_389),
  .S0(ad[5])
);
MUX2 mux_inst_416 (
  .O(mux_o_416),
  .I0(mux_o_390),
  .I1(mux_o_391),
  .S0(ad[5])
);
MUX2 mux_inst_417 (
  .O(mux_o_417),
  .I0(mux_o_392),
  .I1(mux_o_393),
  .S0(ad[5])
);
MUX2 mux_inst_418 (
  .O(mux_o_418),
  .I0(mux_o_394),
  .I1(mux_o_395),
  .S0(ad[5])
);
MUX2 mux_inst_419 (
  .O(mux_o_419),
  .I0(mux_o_396),
  .I1(mux_o_397),
  .S0(ad[5])
);
MUX2 mux_inst_420 (
  .O(mux_o_420),
  .I0(mux_o_398),
  .I1(mux_o_399),
  .S0(ad[5])
);
MUX2 mux_inst_421 (
  .O(mux_o_421),
  .I0(mux_o_400),
  .I1(mux_o_401),
  .S0(ad[5])
);
MUX2 mux_inst_422 (
  .O(mux_o_422),
  .I0(mux_o_402),
  .I1(mux_o_403),
  .S0(ad[5])
);
MUX2 mux_inst_423 (
  .O(mux_o_423),
  .I0(mux_o_404),
  .I1(mux_o_405),
  .S0(ad[5])
);
MUX2 mux_inst_424 (
  .O(mux_o_424),
  .I0(mux_o_406),
  .I1(mux_o_407),
  .S0(ad[5])
);
MUX2 mux_inst_425 (
  .O(mux_o_425),
  .I0(mux_o_408),
  .I1(mux_o_409),
  .S0(ad[5])
);
MUX2 mux_inst_426 (
  .O(mux_o_426),
  .I0(mux_o_410),
  .I1(mux_o_411),
  .S0(ad[6])
);
MUX2 mux_inst_427 (
  .O(mux_o_427),
  .I0(mux_o_412),
  .I1(mux_o_413),
  .S0(ad[6])
);
MUX2 mux_inst_428 (
  .O(mux_o_428),
  .I0(mux_o_414),
  .I1(mux_o_415),
  .S0(ad[6])
);
MUX2 mux_inst_429 (
  .O(mux_o_429),
  .I0(mux_o_416),
  .I1(mux_o_417),
  .S0(ad[6])
);
MUX2 mux_inst_430 (
  .O(mux_o_430),
  .I0(mux_o_418),
  .I1(mux_o_419),
  .S0(ad[6])
);
MUX2 mux_inst_431 (
  .O(mux_o_431),
  .I0(mux_o_420),
  .I1(mux_o_421),
  .S0(ad[6])
);
MUX2 mux_inst_432 (
  .O(mux_o_432),
  .I0(mux_o_422),
  .I1(mux_o_423),
  .S0(ad[6])
);
MUX2 mux_inst_433 (
  .O(mux_o_433),
  .I0(mux_o_424),
  .I1(mux_o_425),
  .S0(ad[6])
);
MUX2 mux_inst_434 (
  .O(mux_o_434),
  .I0(mux_o_426),
  .I1(mux_o_427),
  .S0(ad[7])
);
MUX2 mux_inst_435 (
  .O(mux_o_435),
  .I0(mux_o_428),
  .I1(mux_o_429),
  .S0(ad[7])
);
MUX2 mux_inst_436 (
  .O(mux_o_436),
  .I0(mux_o_430),
  .I1(mux_o_431),
  .S0(ad[7])
);
MUX2 mux_inst_437 (
  .O(mux_o_437),
  .I0(mux_o_432),
  .I1(mux_o_433),
  .S0(ad[7])
);
MUX2 mux_inst_438 (
  .O(mux_o_438),
  .I0(mux_o_434),
  .I1(mux_o_435),
  .S0(ad[8])
);
MUX2 mux_inst_439 (
  .O(mux_o_439),
  .I0(mux_o_436),
  .I1(mux_o_437),
  .S0(ad[8])
);
MUX2 mux_inst_440 (
  .O(dout[6]),
  .I0(mux_o_438),
  .I1(mux_o_439),
  .S0(ad[9])
);
MUX2 mux_inst_441 (
  .O(mux_o_441),
  .I0(rom16_inst_7_dout[7]),
  .I1(rom16_inst_23_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_442 (
  .O(mux_o_442),
  .I0(rom16_inst_39_dout[7]),
  .I1(rom16_inst_55_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_443 (
  .O(mux_o_443),
  .I0(rom16_inst_71_dout[7]),
  .I1(rom16_inst_87_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_444 (
  .O(mux_o_444),
  .I0(rom16_inst_103_dout[7]),
  .I1(rom16_inst_119_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_445 (
  .O(mux_o_445),
  .I0(rom16_inst_135_dout[7]),
  .I1(rom16_inst_151_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_446 (
  .O(mux_o_446),
  .I0(rom16_inst_167_dout[7]),
  .I1(rom16_inst_183_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_447 (
  .O(mux_o_447),
  .I0(rom16_inst_199_dout[7]),
  .I1(rom16_inst_215_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_448 (
  .O(mux_o_448),
  .I0(rom16_inst_231_dout[7]),
  .I1(rom16_inst_247_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_449 (
  .O(mux_o_449),
  .I0(rom16_inst_263_dout[7]),
  .I1(rom16_inst_279_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_450 (
  .O(mux_o_450),
  .I0(rom16_inst_295_dout[7]),
  .I1(rom16_inst_311_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_451 (
  .O(mux_o_451),
  .I0(rom16_inst_327_dout[7]),
  .I1(rom16_inst_343_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_452 (
  .O(mux_o_452),
  .I0(rom16_inst_359_dout[7]),
  .I1(rom16_inst_375_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_453 (
  .O(mux_o_453),
  .I0(rom16_inst_391_dout[7]),
  .I1(rom16_inst_407_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_454 (
  .O(mux_o_454),
  .I0(rom16_inst_423_dout[7]),
  .I1(rom16_inst_439_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_455 (
  .O(mux_o_455),
  .I0(rom16_inst_455_dout[7]),
  .I1(rom16_inst_471_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_456 (
  .O(mux_o_456),
  .I0(rom16_inst_487_dout[7]),
  .I1(rom16_inst_503_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_457 (
  .O(mux_o_457),
  .I0(rom16_inst_519_dout[7]),
  .I1(rom16_inst_535_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_458 (
  .O(mux_o_458),
  .I0(rom16_inst_551_dout[7]),
  .I1(rom16_inst_567_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_459 (
  .O(mux_o_459),
  .I0(rom16_inst_583_dout[7]),
  .I1(rom16_inst_599_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_460 (
  .O(mux_o_460),
  .I0(rom16_inst_615_dout[7]),
  .I1(rom16_inst_631_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_461 (
  .O(mux_o_461),
  .I0(rom16_inst_647_dout[7]),
  .I1(rom16_inst_663_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_462 (
  .O(mux_o_462),
  .I0(rom16_inst_679_dout[7]),
  .I1(rom16_inst_695_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_463 (
  .O(mux_o_463),
  .I0(rom16_inst_711_dout[7]),
  .I1(rom16_inst_727_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_464 (
  .O(mux_o_464),
  .I0(rom16_inst_743_dout[7]),
  .I1(rom16_inst_759_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_465 (
  .O(mux_o_465),
  .I0(rom16_inst_775_dout[7]),
  .I1(rom16_inst_791_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_466 (
  .O(mux_o_466),
  .I0(rom16_inst_807_dout[7]),
  .I1(rom16_inst_823_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_467 (
  .O(mux_o_467),
  .I0(rom16_inst_839_dout[7]),
  .I1(rom16_inst_855_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_468 (
  .O(mux_o_468),
  .I0(rom16_inst_871_dout[7]),
  .I1(rom16_inst_887_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_469 (
  .O(mux_o_469),
  .I0(rom16_inst_903_dout[7]),
  .I1(rom16_inst_919_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_470 (
  .O(mux_o_470),
  .I0(rom16_inst_935_dout[7]),
  .I1(rom16_inst_951_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_471 (
  .O(mux_o_471),
  .I0(rom16_inst_967_dout[7]),
  .I1(rom16_inst_983_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_472 (
  .O(mux_o_472),
  .I0(rom16_inst_999_dout[7]),
  .I1(rom16_inst_1015_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_473 (
  .O(mux_o_473),
  .I0(mux_o_441),
  .I1(mux_o_442),
  .S0(ad[5])
);
MUX2 mux_inst_474 (
  .O(mux_o_474),
  .I0(mux_o_443),
  .I1(mux_o_444),
  .S0(ad[5])
);
MUX2 mux_inst_475 (
  .O(mux_o_475),
  .I0(mux_o_445),
  .I1(mux_o_446),
  .S0(ad[5])
);
MUX2 mux_inst_476 (
  .O(mux_o_476),
  .I0(mux_o_447),
  .I1(mux_o_448),
  .S0(ad[5])
);
MUX2 mux_inst_477 (
  .O(mux_o_477),
  .I0(mux_o_449),
  .I1(mux_o_450),
  .S0(ad[5])
);
MUX2 mux_inst_478 (
  .O(mux_o_478),
  .I0(mux_o_451),
  .I1(mux_o_452),
  .S0(ad[5])
);
MUX2 mux_inst_479 (
  .O(mux_o_479),
  .I0(mux_o_453),
  .I1(mux_o_454),
  .S0(ad[5])
);
MUX2 mux_inst_480 (
  .O(mux_o_480),
  .I0(mux_o_455),
  .I1(mux_o_456),
  .S0(ad[5])
);
MUX2 mux_inst_481 (
  .O(mux_o_481),
  .I0(mux_o_457),
  .I1(mux_o_458),
  .S0(ad[5])
);
MUX2 mux_inst_482 (
  .O(mux_o_482),
  .I0(mux_o_459),
  .I1(mux_o_460),
  .S0(ad[5])
);
MUX2 mux_inst_483 (
  .O(mux_o_483),
  .I0(mux_o_461),
  .I1(mux_o_462),
  .S0(ad[5])
);
MUX2 mux_inst_484 (
  .O(mux_o_484),
  .I0(mux_o_463),
  .I1(mux_o_464),
  .S0(ad[5])
);
MUX2 mux_inst_485 (
  .O(mux_o_485),
  .I0(mux_o_465),
  .I1(mux_o_466),
  .S0(ad[5])
);
MUX2 mux_inst_486 (
  .O(mux_o_486),
  .I0(mux_o_467),
  .I1(mux_o_468),
  .S0(ad[5])
);
MUX2 mux_inst_487 (
  .O(mux_o_487),
  .I0(mux_o_469),
  .I1(mux_o_470),
  .S0(ad[5])
);
MUX2 mux_inst_488 (
  .O(mux_o_488),
  .I0(mux_o_471),
  .I1(mux_o_472),
  .S0(ad[5])
);
MUX2 mux_inst_489 (
  .O(mux_o_489),
  .I0(mux_o_473),
  .I1(mux_o_474),
  .S0(ad[6])
);
MUX2 mux_inst_490 (
  .O(mux_o_490),
  .I0(mux_o_475),
  .I1(mux_o_476),
  .S0(ad[6])
);
MUX2 mux_inst_491 (
  .O(mux_o_491),
  .I0(mux_o_477),
  .I1(mux_o_478),
  .S0(ad[6])
);
MUX2 mux_inst_492 (
  .O(mux_o_492),
  .I0(mux_o_479),
  .I1(mux_o_480),
  .S0(ad[6])
);
MUX2 mux_inst_493 (
  .O(mux_o_493),
  .I0(mux_o_481),
  .I1(mux_o_482),
  .S0(ad[6])
);
MUX2 mux_inst_494 (
  .O(mux_o_494),
  .I0(mux_o_483),
  .I1(mux_o_484),
  .S0(ad[6])
);
MUX2 mux_inst_495 (
  .O(mux_o_495),
  .I0(mux_o_485),
  .I1(mux_o_486),
  .S0(ad[6])
);
MUX2 mux_inst_496 (
  .O(mux_o_496),
  .I0(mux_o_487),
  .I1(mux_o_488),
  .S0(ad[6])
);
MUX2 mux_inst_497 (
  .O(mux_o_497),
  .I0(mux_o_489),
  .I1(mux_o_490),
  .S0(ad[7])
);
MUX2 mux_inst_498 (
  .O(mux_o_498),
  .I0(mux_o_491),
  .I1(mux_o_492),
  .S0(ad[7])
);
MUX2 mux_inst_499 (
  .O(mux_o_499),
  .I0(mux_o_493),
  .I1(mux_o_494),
  .S0(ad[7])
);
MUX2 mux_inst_500 (
  .O(mux_o_500),
  .I0(mux_o_495),
  .I1(mux_o_496),
  .S0(ad[7])
);
MUX2 mux_inst_501 (
  .O(mux_o_501),
  .I0(mux_o_497),
  .I1(mux_o_498),
  .S0(ad[8])
);
MUX2 mux_inst_502 (
  .O(mux_o_502),
  .I0(mux_o_499),
  .I1(mux_o_500),
  .S0(ad[8])
);
MUX2 mux_inst_503 (
  .O(dout[7]),
  .I0(mux_o_501),
  .I1(mux_o_502),
  .S0(ad[9])
);
MUX2 mux_inst_504 (
  .O(mux_o_504),
  .I0(rom16_inst_8_dout[8]),
  .I1(rom16_inst_24_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_505 (
  .O(mux_o_505),
  .I0(rom16_inst_40_dout[8]),
  .I1(rom16_inst_56_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_506 (
  .O(mux_o_506),
  .I0(rom16_inst_72_dout[8]),
  .I1(rom16_inst_88_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_507 (
  .O(mux_o_507),
  .I0(rom16_inst_104_dout[8]),
  .I1(rom16_inst_120_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_508 (
  .O(mux_o_508),
  .I0(rom16_inst_136_dout[8]),
  .I1(rom16_inst_152_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_509 (
  .O(mux_o_509),
  .I0(rom16_inst_168_dout[8]),
  .I1(rom16_inst_184_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_510 (
  .O(mux_o_510),
  .I0(rom16_inst_200_dout[8]),
  .I1(rom16_inst_216_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_511 (
  .O(mux_o_511),
  .I0(rom16_inst_232_dout[8]),
  .I1(rom16_inst_248_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_512 (
  .O(mux_o_512),
  .I0(rom16_inst_264_dout[8]),
  .I1(rom16_inst_280_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_513 (
  .O(mux_o_513),
  .I0(rom16_inst_296_dout[8]),
  .I1(rom16_inst_312_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_514 (
  .O(mux_o_514),
  .I0(rom16_inst_328_dout[8]),
  .I1(rom16_inst_344_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_515 (
  .O(mux_o_515),
  .I0(rom16_inst_360_dout[8]),
  .I1(rom16_inst_376_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_516 (
  .O(mux_o_516),
  .I0(rom16_inst_392_dout[8]),
  .I1(rom16_inst_408_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_517 (
  .O(mux_o_517),
  .I0(rom16_inst_424_dout[8]),
  .I1(rom16_inst_440_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_518 (
  .O(mux_o_518),
  .I0(rom16_inst_456_dout[8]),
  .I1(rom16_inst_472_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_519 (
  .O(mux_o_519),
  .I0(rom16_inst_488_dout[8]),
  .I1(rom16_inst_504_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_520 (
  .O(mux_o_520),
  .I0(rom16_inst_520_dout[8]),
  .I1(rom16_inst_536_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_521 (
  .O(mux_o_521),
  .I0(rom16_inst_552_dout[8]),
  .I1(rom16_inst_568_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_522 (
  .O(mux_o_522),
  .I0(rom16_inst_584_dout[8]),
  .I1(rom16_inst_600_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_523 (
  .O(mux_o_523),
  .I0(rom16_inst_616_dout[8]),
  .I1(rom16_inst_632_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_524 (
  .O(mux_o_524),
  .I0(rom16_inst_648_dout[8]),
  .I1(rom16_inst_664_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_525 (
  .O(mux_o_525),
  .I0(rom16_inst_680_dout[8]),
  .I1(rom16_inst_696_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_526 (
  .O(mux_o_526),
  .I0(rom16_inst_712_dout[8]),
  .I1(rom16_inst_728_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_527 (
  .O(mux_o_527),
  .I0(rom16_inst_744_dout[8]),
  .I1(rom16_inst_760_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_528 (
  .O(mux_o_528),
  .I0(rom16_inst_776_dout[8]),
  .I1(rom16_inst_792_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_529 (
  .O(mux_o_529),
  .I0(rom16_inst_808_dout[8]),
  .I1(rom16_inst_824_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_530 (
  .O(mux_o_530),
  .I0(rom16_inst_840_dout[8]),
  .I1(rom16_inst_856_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_531 (
  .O(mux_o_531),
  .I0(rom16_inst_872_dout[8]),
  .I1(rom16_inst_888_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_532 (
  .O(mux_o_532),
  .I0(rom16_inst_904_dout[8]),
  .I1(rom16_inst_920_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_533 (
  .O(mux_o_533),
  .I0(rom16_inst_936_dout[8]),
  .I1(rom16_inst_952_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_534 (
  .O(mux_o_534),
  .I0(rom16_inst_968_dout[8]),
  .I1(rom16_inst_984_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_535 (
  .O(mux_o_535),
  .I0(rom16_inst_1000_dout[8]),
  .I1(rom16_inst_1016_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_536 (
  .O(mux_o_536),
  .I0(mux_o_504),
  .I1(mux_o_505),
  .S0(ad[5])
);
MUX2 mux_inst_537 (
  .O(mux_o_537),
  .I0(mux_o_506),
  .I1(mux_o_507),
  .S0(ad[5])
);
MUX2 mux_inst_538 (
  .O(mux_o_538),
  .I0(mux_o_508),
  .I1(mux_o_509),
  .S0(ad[5])
);
MUX2 mux_inst_539 (
  .O(mux_o_539),
  .I0(mux_o_510),
  .I1(mux_o_511),
  .S0(ad[5])
);
MUX2 mux_inst_540 (
  .O(mux_o_540),
  .I0(mux_o_512),
  .I1(mux_o_513),
  .S0(ad[5])
);
MUX2 mux_inst_541 (
  .O(mux_o_541),
  .I0(mux_o_514),
  .I1(mux_o_515),
  .S0(ad[5])
);
MUX2 mux_inst_542 (
  .O(mux_o_542),
  .I0(mux_o_516),
  .I1(mux_o_517),
  .S0(ad[5])
);
MUX2 mux_inst_543 (
  .O(mux_o_543),
  .I0(mux_o_518),
  .I1(mux_o_519),
  .S0(ad[5])
);
MUX2 mux_inst_544 (
  .O(mux_o_544),
  .I0(mux_o_520),
  .I1(mux_o_521),
  .S0(ad[5])
);
MUX2 mux_inst_545 (
  .O(mux_o_545),
  .I0(mux_o_522),
  .I1(mux_o_523),
  .S0(ad[5])
);
MUX2 mux_inst_546 (
  .O(mux_o_546),
  .I0(mux_o_524),
  .I1(mux_o_525),
  .S0(ad[5])
);
MUX2 mux_inst_547 (
  .O(mux_o_547),
  .I0(mux_o_526),
  .I1(mux_o_527),
  .S0(ad[5])
);
MUX2 mux_inst_548 (
  .O(mux_o_548),
  .I0(mux_o_528),
  .I1(mux_o_529),
  .S0(ad[5])
);
MUX2 mux_inst_549 (
  .O(mux_o_549),
  .I0(mux_o_530),
  .I1(mux_o_531),
  .S0(ad[5])
);
MUX2 mux_inst_550 (
  .O(mux_o_550),
  .I0(mux_o_532),
  .I1(mux_o_533),
  .S0(ad[5])
);
MUX2 mux_inst_551 (
  .O(mux_o_551),
  .I0(mux_o_534),
  .I1(mux_o_535),
  .S0(ad[5])
);
MUX2 mux_inst_552 (
  .O(mux_o_552),
  .I0(mux_o_536),
  .I1(mux_o_537),
  .S0(ad[6])
);
MUX2 mux_inst_553 (
  .O(mux_o_553),
  .I0(mux_o_538),
  .I1(mux_o_539),
  .S0(ad[6])
);
MUX2 mux_inst_554 (
  .O(mux_o_554),
  .I0(mux_o_540),
  .I1(mux_o_541),
  .S0(ad[6])
);
MUX2 mux_inst_555 (
  .O(mux_o_555),
  .I0(mux_o_542),
  .I1(mux_o_543),
  .S0(ad[6])
);
MUX2 mux_inst_556 (
  .O(mux_o_556),
  .I0(mux_o_544),
  .I1(mux_o_545),
  .S0(ad[6])
);
MUX2 mux_inst_557 (
  .O(mux_o_557),
  .I0(mux_o_546),
  .I1(mux_o_547),
  .S0(ad[6])
);
MUX2 mux_inst_558 (
  .O(mux_o_558),
  .I0(mux_o_548),
  .I1(mux_o_549),
  .S0(ad[6])
);
MUX2 mux_inst_559 (
  .O(mux_o_559),
  .I0(mux_o_550),
  .I1(mux_o_551),
  .S0(ad[6])
);
MUX2 mux_inst_560 (
  .O(mux_o_560),
  .I0(mux_o_552),
  .I1(mux_o_553),
  .S0(ad[7])
);
MUX2 mux_inst_561 (
  .O(mux_o_561),
  .I0(mux_o_554),
  .I1(mux_o_555),
  .S0(ad[7])
);
MUX2 mux_inst_562 (
  .O(mux_o_562),
  .I0(mux_o_556),
  .I1(mux_o_557),
  .S0(ad[7])
);
MUX2 mux_inst_563 (
  .O(mux_o_563),
  .I0(mux_o_558),
  .I1(mux_o_559),
  .S0(ad[7])
);
MUX2 mux_inst_564 (
  .O(mux_o_564),
  .I0(mux_o_560),
  .I1(mux_o_561),
  .S0(ad[8])
);
MUX2 mux_inst_565 (
  .O(mux_o_565),
  .I0(mux_o_562),
  .I1(mux_o_563),
  .S0(ad[8])
);
MUX2 mux_inst_566 (
  .O(dout[8]),
  .I0(mux_o_564),
  .I1(mux_o_565),
  .S0(ad[9])
);
MUX2 mux_inst_567 (
  .O(mux_o_567),
  .I0(rom16_inst_9_dout[9]),
  .I1(rom16_inst_25_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_568 (
  .O(mux_o_568),
  .I0(rom16_inst_41_dout[9]),
  .I1(rom16_inst_57_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_569 (
  .O(mux_o_569),
  .I0(rom16_inst_73_dout[9]),
  .I1(rom16_inst_89_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_570 (
  .O(mux_o_570),
  .I0(rom16_inst_105_dout[9]),
  .I1(rom16_inst_121_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_571 (
  .O(mux_o_571),
  .I0(rom16_inst_137_dout[9]),
  .I1(rom16_inst_153_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_572 (
  .O(mux_o_572),
  .I0(rom16_inst_169_dout[9]),
  .I1(rom16_inst_185_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_573 (
  .O(mux_o_573),
  .I0(rom16_inst_201_dout[9]),
  .I1(rom16_inst_217_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_574 (
  .O(mux_o_574),
  .I0(rom16_inst_233_dout[9]),
  .I1(rom16_inst_249_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_575 (
  .O(mux_o_575),
  .I0(rom16_inst_265_dout[9]),
  .I1(rom16_inst_281_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_576 (
  .O(mux_o_576),
  .I0(rom16_inst_297_dout[9]),
  .I1(rom16_inst_313_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_577 (
  .O(mux_o_577),
  .I0(rom16_inst_329_dout[9]),
  .I1(rom16_inst_345_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_578 (
  .O(mux_o_578),
  .I0(rom16_inst_361_dout[9]),
  .I1(rom16_inst_377_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_579 (
  .O(mux_o_579),
  .I0(rom16_inst_393_dout[9]),
  .I1(rom16_inst_409_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_580 (
  .O(mux_o_580),
  .I0(rom16_inst_425_dout[9]),
  .I1(rom16_inst_441_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_581 (
  .O(mux_o_581),
  .I0(rom16_inst_457_dout[9]),
  .I1(rom16_inst_473_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_582 (
  .O(mux_o_582),
  .I0(rom16_inst_489_dout[9]),
  .I1(rom16_inst_505_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_583 (
  .O(mux_o_583),
  .I0(rom16_inst_521_dout[9]),
  .I1(rom16_inst_537_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_584 (
  .O(mux_o_584),
  .I0(rom16_inst_553_dout[9]),
  .I1(rom16_inst_569_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_585 (
  .O(mux_o_585),
  .I0(rom16_inst_585_dout[9]),
  .I1(rom16_inst_601_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_586 (
  .O(mux_o_586),
  .I0(rom16_inst_617_dout[9]),
  .I1(rom16_inst_633_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_587 (
  .O(mux_o_587),
  .I0(rom16_inst_649_dout[9]),
  .I1(rom16_inst_665_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_588 (
  .O(mux_o_588),
  .I0(rom16_inst_681_dout[9]),
  .I1(rom16_inst_697_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_589 (
  .O(mux_o_589),
  .I0(rom16_inst_713_dout[9]),
  .I1(rom16_inst_729_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_590 (
  .O(mux_o_590),
  .I0(rom16_inst_745_dout[9]),
  .I1(rom16_inst_761_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_591 (
  .O(mux_o_591),
  .I0(rom16_inst_777_dout[9]),
  .I1(rom16_inst_793_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_592 (
  .O(mux_o_592),
  .I0(rom16_inst_809_dout[9]),
  .I1(rom16_inst_825_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_593 (
  .O(mux_o_593),
  .I0(rom16_inst_841_dout[9]),
  .I1(rom16_inst_857_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_594 (
  .O(mux_o_594),
  .I0(rom16_inst_873_dout[9]),
  .I1(rom16_inst_889_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_595 (
  .O(mux_o_595),
  .I0(rom16_inst_905_dout[9]),
  .I1(rom16_inst_921_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_596 (
  .O(mux_o_596),
  .I0(rom16_inst_937_dout[9]),
  .I1(rom16_inst_953_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_597 (
  .O(mux_o_597),
  .I0(rom16_inst_969_dout[9]),
  .I1(rom16_inst_985_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_598 (
  .O(mux_o_598),
  .I0(rom16_inst_1001_dout[9]),
  .I1(rom16_inst_1017_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_599 (
  .O(mux_o_599),
  .I0(mux_o_567),
  .I1(mux_o_568),
  .S0(ad[5])
);
MUX2 mux_inst_600 (
  .O(mux_o_600),
  .I0(mux_o_569),
  .I1(mux_o_570),
  .S0(ad[5])
);
MUX2 mux_inst_601 (
  .O(mux_o_601),
  .I0(mux_o_571),
  .I1(mux_o_572),
  .S0(ad[5])
);
MUX2 mux_inst_602 (
  .O(mux_o_602),
  .I0(mux_o_573),
  .I1(mux_o_574),
  .S0(ad[5])
);
MUX2 mux_inst_603 (
  .O(mux_o_603),
  .I0(mux_o_575),
  .I1(mux_o_576),
  .S0(ad[5])
);
MUX2 mux_inst_604 (
  .O(mux_o_604),
  .I0(mux_o_577),
  .I1(mux_o_578),
  .S0(ad[5])
);
MUX2 mux_inst_605 (
  .O(mux_o_605),
  .I0(mux_o_579),
  .I1(mux_o_580),
  .S0(ad[5])
);
MUX2 mux_inst_606 (
  .O(mux_o_606),
  .I0(mux_o_581),
  .I1(mux_o_582),
  .S0(ad[5])
);
MUX2 mux_inst_607 (
  .O(mux_o_607),
  .I0(mux_o_583),
  .I1(mux_o_584),
  .S0(ad[5])
);
MUX2 mux_inst_608 (
  .O(mux_o_608),
  .I0(mux_o_585),
  .I1(mux_o_586),
  .S0(ad[5])
);
MUX2 mux_inst_609 (
  .O(mux_o_609),
  .I0(mux_o_587),
  .I1(mux_o_588),
  .S0(ad[5])
);
MUX2 mux_inst_610 (
  .O(mux_o_610),
  .I0(mux_o_589),
  .I1(mux_o_590),
  .S0(ad[5])
);
MUX2 mux_inst_611 (
  .O(mux_o_611),
  .I0(mux_o_591),
  .I1(mux_o_592),
  .S0(ad[5])
);
MUX2 mux_inst_612 (
  .O(mux_o_612),
  .I0(mux_o_593),
  .I1(mux_o_594),
  .S0(ad[5])
);
MUX2 mux_inst_613 (
  .O(mux_o_613),
  .I0(mux_o_595),
  .I1(mux_o_596),
  .S0(ad[5])
);
MUX2 mux_inst_614 (
  .O(mux_o_614),
  .I0(mux_o_597),
  .I1(mux_o_598),
  .S0(ad[5])
);
MUX2 mux_inst_615 (
  .O(mux_o_615),
  .I0(mux_o_599),
  .I1(mux_o_600),
  .S0(ad[6])
);
MUX2 mux_inst_616 (
  .O(mux_o_616),
  .I0(mux_o_601),
  .I1(mux_o_602),
  .S0(ad[6])
);
MUX2 mux_inst_617 (
  .O(mux_o_617),
  .I0(mux_o_603),
  .I1(mux_o_604),
  .S0(ad[6])
);
MUX2 mux_inst_618 (
  .O(mux_o_618),
  .I0(mux_o_605),
  .I1(mux_o_606),
  .S0(ad[6])
);
MUX2 mux_inst_619 (
  .O(mux_o_619),
  .I0(mux_o_607),
  .I1(mux_o_608),
  .S0(ad[6])
);
MUX2 mux_inst_620 (
  .O(mux_o_620),
  .I0(mux_o_609),
  .I1(mux_o_610),
  .S0(ad[6])
);
MUX2 mux_inst_621 (
  .O(mux_o_621),
  .I0(mux_o_611),
  .I1(mux_o_612),
  .S0(ad[6])
);
MUX2 mux_inst_622 (
  .O(mux_o_622),
  .I0(mux_o_613),
  .I1(mux_o_614),
  .S0(ad[6])
);
MUX2 mux_inst_623 (
  .O(mux_o_623),
  .I0(mux_o_615),
  .I1(mux_o_616),
  .S0(ad[7])
);
MUX2 mux_inst_624 (
  .O(mux_o_624),
  .I0(mux_o_617),
  .I1(mux_o_618),
  .S0(ad[7])
);
MUX2 mux_inst_625 (
  .O(mux_o_625),
  .I0(mux_o_619),
  .I1(mux_o_620),
  .S0(ad[7])
);
MUX2 mux_inst_626 (
  .O(mux_o_626),
  .I0(mux_o_621),
  .I1(mux_o_622),
  .S0(ad[7])
);
MUX2 mux_inst_627 (
  .O(mux_o_627),
  .I0(mux_o_623),
  .I1(mux_o_624),
  .S0(ad[8])
);
MUX2 mux_inst_628 (
  .O(mux_o_628),
  .I0(mux_o_625),
  .I1(mux_o_626),
  .S0(ad[8])
);
MUX2 mux_inst_629 (
  .O(dout[9]),
  .I0(mux_o_627),
  .I1(mux_o_628),
  .S0(ad[9])
);
MUX2 mux_inst_630 (
  .O(mux_o_630),
  .I0(rom16_inst_10_dout[10]),
  .I1(rom16_inst_26_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_631 (
  .O(mux_o_631),
  .I0(rom16_inst_42_dout[10]),
  .I1(rom16_inst_58_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_632 (
  .O(mux_o_632),
  .I0(rom16_inst_74_dout[10]),
  .I1(rom16_inst_90_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_633 (
  .O(mux_o_633),
  .I0(rom16_inst_106_dout[10]),
  .I1(rom16_inst_122_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_634 (
  .O(mux_o_634),
  .I0(rom16_inst_138_dout[10]),
  .I1(rom16_inst_154_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_635 (
  .O(mux_o_635),
  .I0(rom16_inst_170_dout[10]),
  .I1(rom16_inst_186_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_636 (
  .O(mux_o_636),
  .I0(rom16_inst_202_dout[10]),
  .I1(rom16_inst_218_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_637 (
  .O(mux_o_637),
  .I0(rom16_inst_234_dout[10]),
  .I1(rom16_inst_250_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_638 (
  .O(mux_o_638),
  .I0(rom16_inst_266_dout[10]),
  .I1(rom16_inst_282_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_639 (
  .O(mux_o_639),
  .I0(rom16_inst_298_dout[10]),
  .I1(rom16_inst_314_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_640 (
  .O(mux_o_640),
  .I0(rom16_inst_330_dout[10]),
  .I1(rom16_inst_346_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_641 (
  .O(mux_o_641),
  .I0(rom16_inst_362_dout[10]),
  .I1(rom16_inst_378_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_642 (
  .O(mux_o_642),
  .I0(rom16_inst_394_dout[10]),
  .I1(rom16_inst_410_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_643 (
  .O(mux_o_643),
  .I0(rom16_inst_426_dout[10]),
  .I1(rom16_inst_442_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_644 (
  .O(mux_o_644),
  .I0(rom16_inst_458_dout[10]),
  .I1(rom16_inst_474_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_645 (
  .O(mux_o_645),
  .I0(rom16_inst_490_dout[10]),
  .I1(rom16_inst_506_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_646 (
  .O(mux_o_646),
  .I0(rom16_inst_522_dout[10]),
  .I1(rom16_inst_538_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_647 (
  .O(mux_o_647),
  .I0(rom16_inst_554_dout[10]),
  .I1(rom16_inst_570_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_648 (
  .O(mux_o_648),
  .I0(rom16_inst_586_dout[10]),
  .I1(rom16_inst_602_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_649 (
  .O(mux_o_649),
  .I0(rom16_inst_618_dout[10]),
  .I1(rom16_inst_634_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_650 (
  .O(mux_o_650),
  .I0(rom16_inst_650_dout[10]),
  .I1(rom16_inst_666_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_651 (
  .O(mux_o_651),
  .I0(rom16_inst_682_dout[10]),
  .I1(rom16_inst_698_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_652 (
  .O(mux_o_652),
  .I0(rom16_inst_714_dout[10]),
  .I1(rom16_inst_730_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_653 (
  .O(mux_o_653),
  .I0(rom16_inst_746_dout[10]),
  .I1(rom16_inst_762_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_654 (
  .O(mux_o_654),
  .I0(rom16_inst_778_dout[10]),
  .I1(rom16_inst_794_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_655 (
  .O(mux_o_655),
  .I0(rom16_inst_810_dout[10]),
  .I1(rom16_inst_826_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_656 (
  .O(mux_o_656),
  .I0(rom16_inst_842_dout[10]),
  .I1(rom16_inst_858_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_657 (
  .O(mux_o_657),
  .I0(rom16_inst_874_dout[10]),
  .I1(rom16_inst_890_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_658 (
  .O(mux_o_658),
  .I0(rom16_inst_906_dout[10]),
  .I1(rom16_inst_922_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_659 (
  .O(mux_o_659),
  .I0(rom16_inst_938_dout[10]),
  .I1(rom16_inst_954_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_660 (
  .O(mux_o_660),
  .I0(rom16_inst_970_dout[10]),
  .I1(rom16_inst_986_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_661 (
  .O(mux_o_661),
  .I0(rom16_inst_1002_dout[10]),
  .I1(rom16_inst_1018_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_662 (
  .O(mux_o_662),
  .I0(mux_o_630),
  .I1(mux_o_631),
  .S0(ad[5])
);
MUX2 mux_inst_663 (
  .O(mux_o_663),
  .I0(mux_o_632),
  .I1(mux_o_633),
  .S0(ad[5])
);
MUX2 mux_inst_664 (
  .O(mux_o_664),
  .I0(mux_o_634),
  .I1(mux_o_635),
  .S0(ad[5])
);
MUX2 mux_inst_665 (
  .O(mux_o_665),
  .I0(mux_o_636),
  .I1(mux_o_637),
  .S0(ad[5])
);
MUX2 mux_inst_666 (
  .O(mux_o_666),
  .I0(mux_o_638),
  .I1(mux_o_639),
  .S0(ad[5])
);
MUX2 mux_inst_667 (
  .O(mux_o_667),
  .I0(mux_o_640),
  .I1(mux_o_641),
  .S0(ad[5])
);
MUX2 mux_inst_668 (
  .O(mux_o_668),
  .I0(mux_o_642),
  .I1(mux_o_643),
  .S0(ad[5])
);
MUX2 mux_inst_669 (
  .O(mux_o_669),
  .I0(mux_o_644),
  .I1(mux_o_645),
  .S0(ad[5])
);
MUX2 mux_inst_670 (
  .O(mux_o_670),
  .I0(mux_o_646),
  .I1(mux_o_647),
  .S0(ad[5])
);
MUX2 mux_inst_671 (
  .O(mux_o_671),
  .I0(mux_o_648),
  .I1(mux_o_649),
  .S0(ad[5])
);
MUX2 mux_inst_672 (
  .O(mux_o_672),
  .I0(mux_o_650),
  .I1(mux_o_651),
  .S0(ad[5])
);
MUX2 mux_inst_673 (
  .O(mux_o_673),
  .I0(mux_o_652),
  .I1(mux_o_653),
  .S0(ad[5])
);
MUX2 mux_inst_674 (
  .O(mux_o_674),
  .I0(mux_o_654),
  .I1(mux_o_655),
  .S0(ad[5])
);
MUX2 mux_inst_675 (
  .O(mux_o_675),
  .I0(mux_o_656),
  .I1(mux_o_657),
  .S0(ad[5])
);
MUX2 mux_inst_676 (
  .O(mux_o_676),
  .I0(mux_o_658),
  .I1(mux_o_659),
  .S0(ad[5])
);
MUX2 mux_inst_677 (
  .O(mux_o_677),
  .I0(mux_o_660),
  .I1(mux_o_661),
  .S0(ad[5])
);
MUX2 mux_inst_678 (
  .O(mux_o_678),
  .I0(mux_o_662),
  .I1(mux_o_663),
  .S0(ad[6])
);
MUX2 mux_inst_679 (
  .O(mux_o_679),
  .I0(mux_o_664),
  .I1(mux_o_665),
  .S0(ad[6])
);
MUX2 mux_inst_680 (
  .O(mux_o_680),
  .I0(mux_o_666),
  .I1(mux_o_667),
  .S0(ad[6])
);
MUX2 mux_inst_681 (
  .O(mux_o_681),
  .I0(mux_o_668),
  .I1(mux_o_669),
  .S0(ad[6])
);
MUX2 mux_inst_682 (
  .O(mux_o_682),
  .I0(mux_o_670),
  .I1(mux_o_671),
  .S0(ad[6])
);
MUX2 mux_inst_683 (
  .O(mux_o_683),
  .I0(mux_o_672),
  .I1(mux_o_673),
  .S0(ad[6])
);
MUX2 mux_inst_684 (
  .O(mux_o_684),
  .I0(mux_o_674),
  .I1(mux_o_675),
  .S0(ad[6])
);
MUX2 mux_inst_685 (
  .O(mux_o_685),
  .I0(mux_o_676),
  .I1(mux_o_677),
  .S0(ad[6])
);
MUX2 mux_inst_686 (
  .O(mux_o_686),
  .I0(mux_o_678),
  .I1(mux_o_679),
  .S0(ad[7])
);
MUX2 mux_inst_687 (
  .O(mux_o_687),
  .I0(mux_o_680),
  .I1(mux_o_681),
  .S0(ad[7])
);
MUX2 mux_inst_688 (
  .O(mux_o_688),
  .I0(mux_o_682),
  .I1(mux_o_683),
  .S0(ad[7])
);
MUX2 mux_inst_689 (
  .O(mux_o_689),
  .I0(mux_o_684),
  .I1(mux_o_685),
  .S0(ad[7])
);
MUX2 mux_inst_690 (
  .O(mux_o_690),
  .I0(mux_o_686),
  .I1(mux_o_687),
  .S0(ad[8])
);
MUX2 mux_inst_691 (
  .O(mux_o_691),
  .I0(mux_o_688),
  .I1(mux_o_689),
  .S0(ad[8])
);
MUX2 mux_inst_692 (
  .O(dout[10]),
  .I0(mux_o_690),
  .I1(mux_o_691),
  .S0(ad[9])
);
MUX2 mux_inst_693 (
  .O(mux_o_693),
  .I0(rom16_inst_11_dout[11]),
  .I1(rom16_inst_27_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_694 (
  .O(mux_o_694),
  .I0(rom16_inst_43_dout[11]),
  .I1(rom16_inst_59_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_695 (
  .O(mux_o_695),
  .I0(rom16_inst_75_dout[11]),
  .I1(rom16_inst_91_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_696 (
  .O(mux_o_696),
  .I0(rom16_inst_107_dout[11]),
  .I1(rom16_inst_123_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_697 (
  .O(mux_o_697),
  .I0(rom16_inst_139_dout[11]),
  .I1(rom16_inst_155_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_698 (
  .O(mux_o_698),
  .I0(rom16_inst_171_dout[11]),
  .I1(rom16_inst_187_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_699 (
  .O(mux_o_699),
  .I0(rom16_inst_203_dout[11]),
  .I1(rom16_inst_219_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_700 (
  .O(mux_o_700),
  .I0(rom16_inst_235_dout[11]),
  .I1(rom16_inst_251_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_701 (
  .O(mux_o_701),
  .I0(rom16_inst_267_dout[11]),
  .I1(rom16_inst_283_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_702 (
  .O(mux_o_702),
  .I0(rom16_inst_299_dout[11]),
  .I1(rom16_inst_315_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_703 (
  .O(mux_o_703),
  .I0(rom16_inst_331_dout[11]),
  .I1(rom16_inst_347_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_704 (
  .O(mux_o_704),
  .I0(rom16_inst_363_dout[11]),
  .I1(rom16_inst_379_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_705 (
  .O(mux_o_705),
  .I0(rom16_inst_395_dout[11]),
  .I1(rom16_inst_411_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_706 (
  .O(mux_o_706),
  .I0(rom16_inst_427_dout[11]),
  .I1(rom16_inst_443_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_707 (
  .O(mux_o_707),
  .I0(rom16_inst_459_dout[11]),
  .I1(rom16_inst_475_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_708 (
  .O(mux_o_708),
  .I0(rom16_inst_491_dout[11]),
  .I1(rom16_inst_507_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_709 (
  .O(mux_o_709),
  .I0(rom16_inst_523_dout[11]),
  .I1(rom16_inst_539_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_710 (
  .O(mux_o_710),
  .I0(rom16_inst_555_dout[11]),
  .I1(rom16_inst_571_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_711 (
  .O(mux_o_711),
  .I0(rom16_inst_587_dout[11]),
  .I1(rom16_inst_603_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_712 (
  .O(mux_o_712),
  .I0(rom16_inst_619_dout[11]),
  .I1(rom16_inst_635_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_713 (
  .O(mux_o_713),
  .I0(rom16_inst_651_dout[11]),
  .I1(rom16_inst_667_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_714 (
  .O(mux_o_714),
  .I0(rom16_inst_683_dout[11]),
  .I1(rom16_inst_699_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_715 (
  .O(mux_o_715),
  .I0(rom16_inst_715_dout[11]),
  .I1(rom16_inst_731_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_716 (
  .O(mux_o_716),
  .I0(rom16_inst_747_dout[11]),
  .I1(rom16_inst_763_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_717 (
  .O(mux_o_717),
  .I0(rom16_inst_779_dout[11]),
  .I1(rom16_inst_795_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_718 (
  .O(mux_o_718),
  .I0(rom16_inst_811_dout[11]),
  .I1(rom16_inst_827_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_719 (
  .O(mux_o_719),
  .I0(rom16_inst_843_dout[11]),
  .I1(rom16_inst_859_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_720 (
  .O(mux_o_720),
  .I0(rom16_inst_875_dout[11]),
  .I1(rom16_inst_891_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_721 (
  .O(mux_o_721),
  .I0(rom16_inst_907_dout[11]),
  .I1(rom16_inst_923_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_722 (
  .O(mux_o_722),
  .I0(rom16_inst_939_dout[11]),
  .I1(rom16_inst_955_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_723 (
  .O(mux_o_723),
  .I0(rom16_inst_971_dout[11]),
  .I1(rom16_inst_987_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_724 (
  .O(mux_o_724),
  .I0(rom16_inst_1003_dout[11]),
  .I1(rom16_inst_1019_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_725 (
  .O(mux_o_725),
  .I0(mux_o_693),
  .I1(mux_o_694),
  .S0(ad[5])
);
MUX2 mux_inst_726 (
  .O(mux_o_726),
  .I0(mux_o_695),
  .I1(mux_o_696),
  .S0(ad[5])
);
MUX2 mux_inst_727 (
  .O(mux_o_727),
  .I0(mux_o_697),
  .I1(mux_o_698),
  .S0(ad[5])
);
MUX2 mux_inst_728 (
  .O(mux_o_728),
  .I0(mux_o_699),
  .I1(mux_o_700),
  .S0(ad[5])
);
MUX2 mux_inst_729 (
  .O(mux_o_729),
  .I0(mux_o_701),
  .I1(mux_o_702),
  .S0(ad[5])
);
MUX2 mux_inst_730 (
  .O(mux_o_730),
  .I0(mux_o_703),
  .I1(mux_o_704),
  .S0(ad[5])
);
MUX2 mux_inst_731 (
  .O(mux_o_731),
  .I0(mux_o_705),
  .I1(mux_o_706),
  .S0(ad[5])
);
MUX2 mux_inst_732 (
  .O(mux_o_732),
  .I0(mux_o_707),
  .I1(mux_o_708),
  .S0(ad[5])
);
MUX2 mux_inst_733 (
  .O(mux_o_733),
  .I0(mux_o_709),
  .I1(mux_o_710),
  .S0(ad[5])
);
MUX2 mux_inst_734 (
  .O(mux_o_734),
  .I0(mux_o_711),
  .I1(mux_o_712),
  .S0(ad[5])
);
MUX2 mux_inst_735 (
  .O(mux_o_735),
  .I0(mux_o_713),
  .I1(mux_o_714),
  .S0(ad[5])
);
MUX2 mux_inst_736 (
  .O(mux_o_736),
  .I0(mux_o_715),
  .I1(mux_o_716),
  .S0(ad[5])
);
MUX2 mux_inst_737 (
  .O(mux_o_737),
  .I0(mux_o_717),
  .I1(mux_o_718),
  .S0(ad[5])
);
MUX2 mux_inst_738 (
  .O(mux_o_738),
  .I0(mux_o_719),
  .I1(mux_o_720),
  .S0(ad[5])
);
MUX2 mux_inst_739 (
  .O(mux_o_739),
  .I0(mux_o_721),
  .I1(mux_o_722),
  .S0(ad[5])
);
MUX2 mux_inst_740 (
  .O(mux_o_740),
  .I0(mux_o_723),
  .I1(mux_o_724),
  .S0(ad[5])
);
MUX2 mux_inst_741 (
  .O(mux_o_741),
  .I0(mux_o_725),
  .I1(mux_o_726),
  .S0(ad[6])
);
MUX2 mux_inst_742 (
  .O(mux_o_742),
  .I0(mux_o_727),
  .I1(mux_o_728),
  .S0(ad[6])
);
MUX2 mux_inst_743 (
  .O(mux_o_743),
  .I0(mux_o_729),
  .I1(mux_o_730),
  .S0(ad[6])
);
MUX2 mux_inst_744 (
  .O(mux_o_744),
  .I0(mux_o_731),
  .I1(mux_o_732),
  .S0(ad[6])
);
MUX2 mux_inst_745 (
  .O(mux_o_745),
  .I0(mux_o_733),
  .I1(mux_o_734),
  .S0(ad[6])
);
MUX2 mux_inst_746 (
  .O(mux_o_746),
  .I0(mux_o_735),
  .I1(mux_o_736),
  .S0(ad[6])
);
MUX2 mux_inst_747 (
  .O(mux_o_747),
  .I0(mux_o_737),
  .I1(mux_o_738),
  .S0(ad[6])
);
MUX2 mux_inst_748 (
  .O(mux_o_748),
  .I0(mux_o_739),
  .I1(mux_o_740),
  .S0(ad[6])
);
MUX2 mux_inst_749 (
  .O(mux_o_749),
  .I0(mux_o_741),
  .I1(mux_o_742),
  .S0(ad[7])
);
MUX2 mux_inst_750 (
  .O(mux_o_750),
  .I0(mux_o_743),
  .I1(mux_o_744),
  .S0(ad[7])
);
MUX2 mux_inst_751 (
  .O(mux_o_751),
  .I0(mux_o_745),
  .I1(mux_o_746),
  .S0(ad[7])
);
MUX2 mux_inst_752 (
  .O(mux_o_752),
  .I0(mux_o_747),
  .I1(mux_o_748),
  .S0(ad[7])
);
MUX2 mux_inst_753 (
  .O(mux_o_753),
  .I0(mux_o_749),
  .I1(mux_o_750),
  .S0(ad[8])
);
MUX2 mux_inst_754 (
  .O(mux_o_754),
  .I0(mux_o_751),
  .I1(mux_o_752),
  .S0(ad[8])
);
MUX2 mux_inst_755 (
  .O(dout[11]),
  .I0(mux_o_753),
  .I1(mux_o_754),
  .S0(ad[9])
);
MUX2 mux_inst_756 (
  .O(mux_o_756),
  .I0(rom16_inst_12_dout[12]),
  .I1(rom16_inst_28_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_757 (
  .O(mux_o_757),
  .I0(rom16_inst_44_dout[12]),
  .I1(rom16_inst_60_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_758 (
  .O(mux_o_758),
  .I0(rom16_inst_76_dout[12]),
  .I1(rom16_inst_92_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_759 (
  .O(mux_o_759),
  .I0(rom16_inst_108_dout[12]),
  .I1(rom16_inst_124_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_760 (
  .O(mux_o_760),
  .I0(rom16_inst_140_dout[12]),
  .I1(rom16_inst_156_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_761 (
  .O(mux_o_761),
  .I0(rom16_inst_172_dout[12]),
  .I1(rom16_inst_188_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_762 (
  .O(mux_o_762),
  .I0(rom16_inst_204_dout[12]),
  .I1(rom16_inst_220_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_763 (
  .O(mux_o_763),
  .I0(rom16_inst_236_dout[12]),
  .I1(rom16_inst_252_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_764 (
  .O(mux_o_764),
  .I0(rom16_inst_268_dout[12]),
  .I1(rom16_inst_284_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_765 (
  .O(mux_o_765),
  .I0(rom16_inst_300_dout[12]),
  .I1(rom16_inst_316_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_766 (
  .O(mux_o_766),
  .I0(rom16_inst_332_dout[12]),
  .I1(rom16_inst_348_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_767 (
  .O(mux_o_767),
  .I0(rom16_inst_364_dout[12]),
  .I1(rom16_inst_380_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_768 (
  .O(mux_o_768),
  .I0(rom16_inst_396_dout[12]),
  .I1(rom16_inst_412_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_769 (
  .O(mux_o_769),
  .I0(rom16_inst_428_dout[12]),
  .I1(rom16_inst_444_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_770 (
  .O(mux_o_770),
  .I0(rom16_inst_460_dout[12]),
  .I1(rom16_inst_476_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_771 (
  .O(mux_o_771),
  .I0(rom16_inst_492_dout[12]),
  .I1(rom16_inst_508_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_772 (
  .O(mux_o_772),
  .I0(rom16_inst_524_dout[12]),
  .I1(rom16_inst_540_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_773 (
  .O(mux_o_773),
  .I0(rom16_inst_556_dout[12]),
  .I1(rom16_inst_572_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_774 (
  .O(mux_o_774),
  .I0(rom16_inst_588_dout[12]),
  .I1(rom16_inst_604_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_775 (
  .O(mux_o_775),
  .I0(rom16_inst_620_dout[12]),
  .I1(rom16_inst_636_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_776 (
  .O(mux_o_776),
  .I0(rom16_inst_652_dout[12]),
  .I1(rom16_inst_668_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_777 (
  .O(mux_o_777),
  .I0(rom16_inst_684_dout[12]),
  .I1(rom16_inst_700_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_778 (
  .O(mux_o_778),
  .I0(rom16_inst_716_dout[12]),
  .I1(rom16_inst_732_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_779 (
  .O(mux_o_779),
  .I0(rom16_inst_748_dout[12]),
  .I1(rom16_inst_764_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_780 (
  .O(mux_o_780),
  .I0(rom16_inst_780_dout[12]),
  .I1(rom16_inst_796_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_781 (
  .O(mux_o_781),
  .I0(rom16_inst_812_dout[12]),
  .I1(rom16_inst_828_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_782 (
  .O(mux_o_782),
  .I0(rom16_inst_844_dout[12]),
  .I1(rom16_inst_860_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_783 (
  .O(mux_o_783),
  .I0(rom16_inst_876_dout[12]),
  .I1(rom16_inst_892_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_784 (
  .O(mux_o_784),
  .I0(rom16_inst_908_dout[12]),
  .I1(rom16_inst_924_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_785 (
  .O(mux_o_785),
  .I0(rom16_inst_940_dout[12]),
  .I1(rom16_inst_956_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_786 (
  .O(mux_o_786),
  .I0(rom16_inst_972_dout[12]),
  .I1(rom16_inst_988_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_787 (
  .O(mux_o_787),
  .I0(rom16_inst_1004_dout[12]),
  .I1(rom16_inst_1020_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_788 (
  .O(mux_o_788),
  .I0(mux_o_756),
  .I1(mux_o_757),
  .S0(ad[5])
);
MUX2 mux_inst_789 (
  .O(mux_o_789),
  .I0(mux_o_758),
  .I1(mux_o_759),
  .S0(ad[5])
);
MUX2 mux_inst_790 (
  .O(mux_o_790),
  .I0(mux_o_760),
  .I1(mux_o_761),
  .S0(ad[5])
);
MUX2 mux_inst_791 (
  .O(mux_o_791),
  .I0(mux_o_762),
  .I1(mux_o_763),
  .S0(ad[5])
);
MUX2 mux_inst_792 (
  .O(mux_o_792),
  .I0(mux_o_764),
  .I1(mux_o_765),
  .S0(ad[5])
);
MUX2 mux_inst_793 (
  .O(mux_o_793),
  .I0(mux_o_766),
  .I1(mux_o_767),
  .S0(ad[5])
);
MUX2 mux_inst_794 (
  .O(mux_o_794),
  .I0(mux_o_768),
  .I1(mux_o_769),
  .S0(ad[5])
);
MUX2 mux_inst_795 (
  .O(mux_o_795),
  .I0(mux_o_770),
  .I1(mux_o_771),
  .S0(ad[5])
);
MUX2 mux_inst_796 (
  .O(mux_o_796),
  .I0(mux_o_772),
  .I1(mux_o_773),
  .S0(ad[5])
);
MUX2 mux_inst_797 (
  .O(mux_o_797),
  .I0(mux_o_774),
  .I1(mux_o_775),
  .S0(ad[5])
);
MUX2 mux_inst_798 (
  .O(mux_o_798),
  .I0(mux_o_776),
  .I1(mux_o_777),
  .S0(ad[5])
);
MUX2 mux_inst_799 (
  .O(mux_o_799),
  .I0(mux_o_778),
  .I1(mux_o_779),
  .S0(ad[5])
);
MUX2 mux_inst_800 (
  .O(mux_o_800),
  .I0(mux_o_780),
  .I1(mux_o_781),
  .S0(ad[5])
);
MUX2 mux_inst_801 (
  .O(mux_o_801),
  .I0(mux_o_782),
  .I1(mux_o_783),
  .S0(ad[5])
);
MUX2 mux_inst_802 (
  .O(mux_o_802),
  .I0(mux_o_784),
  .I1(mux_o_785),
  .S0(ad[5])
);
MUX2 mux_inst_803 (
  .O(mux_o_803),
  .I0(mux_o_786),
  .I1(mux_o_787),
  .S0(ad[5])
);
MUX2 mux_inst_804 (
  .O(mux_o_804),
  .I0(mux_o_788),
  .I1(mux_o_789),
  .S0(ad[6])
);
MUX2 mux_inst_805 (
  .O(mux_o_805),
  .I0(mux_o_790),
  .I1(mux_o_791),
  .S0(ad[6])
);
MUX2 mux_inst_806 (
  .O(mux_o_806),
  .I0(mux_o_792),
  .I1(mux_o_793),
  .S0(ad[6])
);
MUX2 mux_inst_807 (
  .O(mux_o_807),
  .I0(mux_o_794),
  .I1(mux_o_795),
  .S0(ad[6])
);
MUX2 mux_inst_808 (
  .O(mux_o_808),
  .I0(mux_o_796),
  .I1(mux_o_797),
  .S0(ad[6])
);
MUX2 mux_inst_809 (
  .O(mux_o_809),
  .I0(mux_o_798),
  .I1(mux_o_799),
  .S0(ad[6])
);
MUX2 mux_inst_810 (
  .O(mux_o_810),
  .I0(mux_o_800),
  .I1(mux_o_801),
  .S0(ad[6])
);
MUX2 mux_inst_811 (
  .O(mux_o_811),
  .I0(mux_o_802),
  .I1(mux_o_803),
  .S0(ad[6])
);
MUX2 mux_inst_812 (
  .O(mux_o_812),
  .I0(mux_o_804),
  .I1(mux_o_805),
  .S0(ad[7])
);
MUX2 mux_inst_813 (
  .O(mux_o_813),
  .I0(mux_o_806),
  .I1(mux_o_807),
  .S0(ad[7])
);
MUX2 mux_inst_814 (
  .O(mux_o_814),
  .I0(mux_o_808),
  .I1(mux_o_809),
  .S0(ad[7])
);
MUX2 mux_inst_815 (
  .O(mux_o_815),
  .I0(mux_o_810),
  .I1(mux_o_811),
  .S0(ad[7])
);
MUX2 mux_inst_816 (
  .O(mux_o_816),
  .I0(mux_o_812),
  .I1(mux_o_813),
  .S0(ad[8])
);
MUX2 mux_inst_817 (
  .O(mux_o_817),
  .I0(mux_o_814),
  .I1(mux_o_815),
  .S0(ad[8])
);
MUX2 mux_inst_818 (
  .O(dout[12]),
  .I0(mux_o_816),
  .I1(mux_o_817),
  .S0(ad[9])
);
MUX2 mux_inst_819 (
  .O(mux_o_819),
  .I0(rom16_inst_13_dout[13]),
  .I1(rom16_inst_29_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_820 (
  .O(mux_o_820),
  .I0(rom16_inst_45_dout[13]),
  .I1(rom16_inst_61_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_821 (
  .O(mux_o_821),
  .I0(rom16_inst_77_dout[13]),
  .I1(rom16_inst_93_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_822 (
  .O(mux_o_822),
  .I0(rom16_inst_109_dout[13]),
  .I1(rom16_inst_125_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_823 (
  .O(mux_o_823),
  .I0(rom16_inst_141_dout[13]),
  .I1(rom16_inst_157_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_824 (
  .O(mux_o_824),
  .I0(rom16_inst_173_dout[13]),
  .I1(rom16_inst_189_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_825 (
  .O(mux_o_825),
  .I0(rom16_inst_205_dout[13]),
  .I1(rom16_inst_221_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_826 (
  .O(mux_o_826),
  .I0(rom16_inst_237_dout[13]),
  .I1(rom16_inst_253_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_827 (
  .O(mux_o_827),
  .I0(rom16_inst_269_dout[13]),
  .I1(rom16_inst_285_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_828 (
  .O(mux_o_828),
  .I0(rom16_inst_301_dout[13]),
  .I1(rom16_inst_317_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_829 (
  .O(mux_o_829),
  .I0(rom16_inst_333_dout[13]),
  .I1(rom16_inst_349_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_830 (
  .O(mux_o_830),
  .I0(rom16_inst_365_dout[13]),
  .I1(rom16_inst_381_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_831 (
  .O(mux_o_831),
  .I0(rom16_inst_397_dout[13]),
  .I1(rom16_inst_413_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_832 (
  .O(mux_o_832),
  .I0(rom16_inst_429_dout[13]),
  .I1(rom16_inst_445_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_833 (
  .O(mux_o_833),
  .I0(rom16_inst_461_dout[13]),
  .I1(rom16_inst_477_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_834 (
  .O(mux_o_834),
  .I0(rom16_inst_493_dout[13]),
  .I1(rom16_inst_509_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_835 (
  .O(mux_o_835),
  .I0(rom16_inst_525_dout[13]),
  .I1(rom16_inst_541_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_836 (
  .O(mux_o_836),
  .I0(rom16_inst_557_dout[13]),
  .I1(rom16_inst_573_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_837 (
  .O(mux_o_837),
  .I0(rom16_inst_589_dout[13]),
  .I1(rom16_inst_605_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_838 (
  .O(mux_o_838),
  .I0(rom16_inst_621_dout[13]),
  .I1(rom16_inst_637_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_839 (
  .O(mux_o_839),
  .I0(rom16_inst_653_dout[13]),
  .I1(rom16_inst_669_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_840 (
  .O(mux_o_840),
  .I0(rom16_inst_685_dout[13]),
  .I1(rom16_inst_701_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_841 (
  .O(mux_o_841),
  .I0(rom16_inst_717_dout[13]),
  .I1(rom16_inst_733_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_842 (
  .O(mux_o_842),
  .I0(rom16_inst_749_dout[13]),
  .I1(rom16_inst_765_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_843 (
  .O(mux_o_843),
  .I0(rom16_inst_781_dout[13]),
  .I1(rom16_inst_797_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_844 (
  .O(mux_o_844),
  .I0(rom16_inst_813_dout[13]),
  .I1(rom16_inst_829_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_845 (
  .O(mux_o_845),
  .I0(rom16_inst_845_dout[13]),
  .I1(rom16_inst_861_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_846 (
  .O(mux_o_846),
  .I0(rom16_inst_877_dout[13]),
  .I1(rom16_inst_893_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_847 (
  .O(mux_o_847),
  .I0(rom16_inst_909_dout[13]),
  .I1(rom16_inst_925_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_848 (
  .O(mux_o_848),
  .I0(rom16_inst_941_dout[13]),
  .I1(rom16_inst_957_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_849 (
  .O(mux_o_849),
  .I0(rom16_inst_973_dout[13]),
  .I1(rom16_inst_989_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_850 (
  .O(mux_o_850),
  .I0(rom16_inst_1005_dout[13]),
  .I1(rom16_inst_1021_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_851 (
  .O(mux_o_851),
  .I0(mux_o_819),
  .I1(mux_o_820),
  .S0(ad[5])
);
MUX2 mux_inst_852 (
  .O(mux_o_852),
  .I0(mux_o_821),
  .I1(mux_o_822),
  .S0(ad[5])
);
MUX2 mux_inst_853 (
  .O(mux_o_853),
  .I0(mux_o_823),
  .I1(mux_o_824),
  .S0(ad[5])
);
MUX2 mux_inst_854 (
  .O(mux_o_854),
  .I0(mux_o_825),
  .I1(mux_o_826),
  .S0(ad[5])
);
MUX2 mux_inst_855 (
  .O(mux_o_855),
  .I0(mux_o_827),
  .I1(mux_o_828),
  .S0(ad[5])
);
MUX2 mux_inst_856 (
  .O(mux_o_856),
  .I0(mux_o_829),
  .I1(mux_o_830),
  .S0(ad[5])
);
MUX2 mux_inst_857 (
  .O(mux_o_857),
  .I0(mux_o_831),
  .I1(mux_o_832),
  .S0(ad[5])
);
MUX2 mux_inst_858 (
  .O(mux_o_858),
  .I0(mux_o_833),
  .I1(mux_o_834),
  .S0(ad[5])
);
MUX2 mux_inst_859 (
  .O(mux_o_859),
  .I0(mux_o_835),
  .I1(mux_o_836),
  .S0(ad[5])
);
MUX2 mux_inst_860 (
  .O(mux_o_860),
  .I0(mux_o_837),
  .I1(mux_o_838),
  .S0(ad[5])
);
MUX2 mux_inst_861 (
  .O(mux_o_861),
  .I0(mux_o_839),
  .I1(mux_o_840),
  .S0(ad[5])
);
MUX2 mux_inst_862 (
  .O(mux_o_862),
  .I0(mux_o_841),
  .I1(mux_o_842),
  .S0(ad[5])
);
MUX2 mux_inst_863 (
  .O(mux_o_863),
  .I0(mux_o_843),
  .I1(mux_o_844),
  .S0(ad[5])
);
MUX2 mux_inst_864 (
  .O(mux_o_864),
  .I0(mux_o_845),
  .I1(mux_o_846),
  .S0(ad[5])
);
MUX2 mux_inst_865 (
  .O(mux_o_865),
  .I0(mux_o_847),
  .I1(mux_o_848),
  .S0(ad[5])
);
MUX2 mux_inst_866 (
  .O(mux_o_866),
  .I0(mux_o_849),
  .I1(mux_o_850),
  .S0(ad[5])
);
MUX2 mux_inst_867 (
  .O(mux_o_867),
  .I0(mux_o_851),
  .I1(mux_o_852),
  .S0(ad[6])
);
MUX2 mux_inst_868 (
  .O(mux_o_868),
  .I0(mux_o_853),
  .I1(mux_o_854),
  .S0(ad[6])
);
MUX2 mux_inst_869 (
  .O(mux_o_869),
  .I0(mux_o_855),
  .I1(mux_o_856),
  .S0(ad[6])
);
MUX2 mux_inst_870 (
  .O(mux_o_870),
  .I0(mux_o_857),
  .I1(mux_o_858),
  .S0(ad[6])
);
MUX2 mux_inst_871 (
  .O(mux_o_871),
  .I0(mux_o_859),
  .I1(mux_o_860),
  .S0(ad[6])
);
MUX2 mux_inst_872 (
  .O(mux_o_872),
  .I0(mux_o_861),
  .I1(mux_o_862),
  .S0(ad[6])
);
MUX2 mux_inst_873 (
  .O(mux_o_873),
  .I0(mux_o_863),
  .I1(mux_o_864),
  .S0(ad[6])
);
MUX2 mux_inst_874 (
  .O(mux_o_874),
  .I0(mux_o_865),
  .I1(mux_o_866),
  .S0(ad[6])
);
MUX2 mux_inst_875 (
  .O(mux_o_875),
  .I0(mux_o_867),
  .I1(mux_o_868),
  .S0(ad[7])
);
MUX2 mux_inst_876 (
  .O(mux_o_876),
  .I0(mux_o_869),
  .I1(mux_o_870),
  .S0(ad[7])
);
MUX2 mux_inst_877 (
  .O(mux_o_877),
  .I0(mux_o_871),
  .I1(mux_o_872),
  .S0(ad[7])
);
MUX2 mux_inst_878 (
  .O(mux_o_878),
  .I0(mux_o_873),
  .I1(mux_o_874),
  .S0(ad[7])
);
MUX2 mux_inst_879 (
  .O(mux_o_879),
  .I0(mux_o_875),
  .I1(mux_o_876),
  .S0(ad[8])
);
MUX2 mux_inst_880 (
  .O(mux_o_880),
  .I0(mux_o_877),
  .I1(mux_o_878),
  .S0(ad[8])
);
MUX2 mux_inst_881 (
  .O(dout[13]),
  .I0(mux_o_879),
  .I1(mux_o_880),
  .S0(ad[9])
);
MUX2 mux_inst_882 (
  .O(mux_o_882),
  .I0(rom16_inst_14_dout[14]),
  .I1(rom16_inst_30_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_883 (
  .O(mux_o_883),
  .I0(rom16_inst_46_dout[14]),
  .I1(rom16_inst_62_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_884 (
  .O(mux_o_884),
  .I0(rom16_inst_78_dout[14]),
  .I1(rom16_inst_94_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_885 (
  .O(mux_o_885),
  .I0(rom16_inst_110_dout[14]),
  .I1(rom16_inst_126_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_886 (
  .O(mux_o_886),
  .I0(rom16_inst_142_dout[14]),
  .I1(rom16_inst_158_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_887 (
  .O(mux_o_887),
  .I0(rom16_inst_174_dout[14]),
  .I1(rom16_inst_190_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_888 (
  .O(mux_o_888),
  .I0(rom16_inst_206_dout[14]),
  .I1(rom16_inst_222_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_889 (
  .O(mux_o_889),
  .I0(rom16_inst_238_dout[14]),
  .I1(rom16_inst_254_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_890 (
  .O(mux_o_890),
  .I0(rom16_inst_270_dout[14]),
  .I1(rom16_inst_286_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_891 (
  .O(mux_o_891),
  .I0(rom16_inst_302_dout[14]),
  .I1(rom16_inst_318_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_892 (
  .O(mux_o_892),
  .I0(rom16_inst_334_dout[14]),
  .I1(rom16_inst_350_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_893 (
  .O(mux_o_893),
  .I0(rom16_inst_366_dout[14]),
  .I1(rom16_inst_382_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_894 (
  .O(mux_o_894),
  .I0(rom16_inst_398_dout[14]),
  .I1(rom16_inst_414_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_895 (
  .O(mux_o_895),
  .I0(rom16_inst_430_dout[14]),
  .I1(rom16_inst_446_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_896 (
  .O(mux_o_896),
  .I0(rom16_inst_462_dout[14]),
  .I1(rom16_inst_478_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_897 (
  .O(mux_o_897),
  .I0(rom16_inst_494_dout[14]),
  .I1(rom16_inst_510_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_898 (
  .O(mux_o_898),
  .I0(rom16_inst_526_dout[14]),
  .I1(rom16_inst_542_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_899 (
  .O(mux_o_899),
  .I0(rom16_inst_558_dout[14]),
  .I1(rom16_inst_574_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_900 (
  .O(mux_o_900),
  .I0(rom16_inst_590_dout[14]),
  .I1(rom16_inst_606_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_901 (
  .O(mux_o_901),
  .I0(rom16_inst_622_dout[14]),
  .I1(rom16_inst_638_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_902 (
  .O(mux_o_902),
  .I0(rom16_inst_654_dout[14]),
  .I1(rom16_inst_670_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_903 (
  .O(mux_o_903),
  .I0(rom16_inst_686_dout[14]),
  .I1(rom16_inst_702_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_904 (
  .O(mux_o_904),
  .I0(rom16_inst_718_dout[14]),
  .I1(rom16_inst_734_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_905 (
  .O(mux_o_905),
  .I0(rom16_inst_750_dout[14]),
  .I1(rom16_inst_766_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_906 (
  .O(mux_o_906),
  .I0(rom16_inst_782_dout[14]),
  .I1(rom16_inst_798_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_907 (
  .O(mux_o_907),
  .I0(rom16_inst_814_dout[14]),
  .I1(rom16_inst_830_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_908 (
  .O(mux_o_908),
  .I0(rom16_inst_846_dout[14]),
  .I1(rom16_inst_862_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_909 (
  .O(mux_o_909),
  .I0(rom16_inst_878_dout[14]),
  .I1(rom16_inst_894_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_910 (
  .O(mux_o_910),
  .I0(rom16_inst_910_dout[14]),
  .I1(rom16_inst_926_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_911 (
  .O(mux_o_911),
  .I0(rom16_inst_942_dout[14]),
  .I1(rom16_inst_958_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_912 (
  .O(mux_o_912),
  .I0(rom16_inst_974_dout[14]),
  .I1(rom16_inst_990_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_913 (
  .O(mux_o_913),
  .I0(rom16_inst_1006_dout[14]),
  .I1(rom16_inst_1022_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_914 (
  .O(mux_o_914),
  .I0(mux_o_882),
  .I1(mux_o_883),
  .S0(ad[5])
);
MUX2 mux_inst_915 (
  .O(mux_o_915),
  .I0(mux_o_884),
  .I1(mux_o_885),
  .S0(ad[5])
);
MUX2 mux_inst_916 (
  .O(mux_o_916),
  .I0(mux_o_886),
  .I1(mux_o_887),
  .S0(ad[5])
);
MUX2 mux_inst_917 (
  .O(mux_o_917),
  .I0(mux_o_888),
  .I1(mux_o_889),
  .S0(ad[5])
);
MUX2 mux_inst_918 (
  .O(mux_o_918),
  .I0(mux_o_890),
  .I1(mux_o_891),
  .S0(ad[5])
);
MUX2 mux_inst_919 (
  .O(mux_o_919),
  .I0(mux_o_892),
  .I1(mux_o_893),
  .S0(ad[5])
);
MUX2 mux_inst_920 (
  .O(mux_o_920),
  .I0(mux_o_894),
  .I1(mux_o_895),
  .S0(ad[5])
);
MUX2 mux_inst_921 (
  .O(mux_o_921),
  .I0(mux_o_896),
  .I1(mux_o_897),
  .S0(ad[5])
);
MUX2 mux_inst_922 (
  .O(mux_o_922),
  .I0(mux_o_898),
  .I1(mux_o_899),
  .S0(ad[5])
);
MUX2 mux_inst_923 (
  .O(mux_o_923),
  .I0(mux_o_900),
  .I1(mux_o_901),
  .S0(ad[5])
);
MUX2 mux_inst_924 (
  .O(mux_o_924),
  .I0(mux_o_902),
  .I1(mux_o_903),
  .S0(ad[5])
);
MUX2 mux_inst_925 (
  .O(mux_o_925),
  .I0(mux_o_904),
  .I1(mux_o_905),
  .S0(ad[5])
);
MUX2 mux_inst_926 (
  .O(mux_o_926),
  .I0(mux_o_906),
  .I1(mux_o_907),
  .S0(ad[5])
);
MUX2 mux_inst_927 (
  .O(mux_o_927),
  .I0(mux_o_908),
  .I1(mux_o_909),
  .S0(ad[5])
);
MUX2 mux_inst_928 (
  .O(mux_o_928),
  .I0(mux_o_910),
  .I1(mux_o_911),
  .S0(ad[5])
);
MUX2 mux_inst_929 (
  .O(mux_o_929),
  .I0(mux_o_912),
  .I1(mux_o_913),
  .S0(ad[5])
);
MUX2 mux_inst_930 (
  .O(mux_o_930),
  .I0(mux_o_914),
  .I1(mux_o_915),
  .S0(ad[6])
);
MUX2 mux_inst_931 (
  .O(mux_o_931),
  .I0(mux_o_916),
  .I1(mux_o_917),
  .S0(ad[6])
);
MUX2 mux_inst_932 (
  .O(mux_o_932),
  .I0(mux_o_918),
  .I1(mux_o_919),
  .S0(ad[6])
);
MUX2 mux_inst_933 (
  .O(mux_o_933),
  .I0(mux_o_920),
  .I1(mux_o_921),
  .S0(ad[6])
);
MUX2 mux_inst_934 (
  .O(mux_o_934),
  .I0(mux_o_922),
  .I1(mux_o_923),
  .S0(ad[6])
);
MUX2 mux_inst_935 (
  .O(mux_o_935),
  .I0(mux_o_924),
  .I1(mux_o_925),
  .S0(ad[6])
);
MUX2 mux_inst_936 (
  .O(mux_o_936),
  .I0(mux_o_926),
  .I1(mux_o_927),
  .S0(ad[6])
);
MUX2 mux_inst_937 (
  .O(mux_o_937),
  .I0(mux_o_928),
  .I1(mux_o_929),
  .S0(ad[6])
);
MUX2 mux_inst_938 (
  .O(mux_o_938),
  .I0(mux_o_930),
  .I1(mux_o_931),
  .S0(ad[7])
);
MUX2 mux_inst_939 (
  .O(mux_o_939),
  .I0(mux_o_932),
  .I1(mux_o_933),
  .S0(ad[7])
);
MUX2 mux_inst_940 (
  .O(mux_o_940),
  .I0(mux_o_934),
  .I1(mux_o_935),
  .S0(ad[7])
);
MUX2 mux_inst_941 (
  .O(mux_o_941),
  .I0(mux_o_936),
  .I1(mux_o_937),
  .S0(ad[7])
);
MUX2 mux_inst_942 (
  .O(mux_o_942),
  .I0(mux_o_938),
  .I1(mux_o_939),
  .S0(ad[8])
);
MUX2 mux_inst_943 (
  .O(mux_o_943),
  .I0(mux_o_940),
  .I1(mux_o_941),
  .S0(ad[8])
);
MUX2 mux_inst_944 (
  .O(dout[14]),
  .I0(mux_o_942),
  .I1(mux_o_943),
  .S0(ad[9])
);
MUX2 mux_inst_945 (
  .O(mux_o_945),
  .I0(rom16_inst_15_dout[15]),
  .I1(rom16_inst_31_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_946 (
  .O(mux_o_946),
  .I0(rom16_inst_47_dout[15]),
  .I1(rom16_inst_63_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_947 (
  .O(mux_o_947),
  .I0(rom16_inst_79_dout[15]),
  .I1(rom16_inst_95_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_948 (
  .O(mux_o_948),
  .I0(rom16_inst_111_dout[15]),
  .I1(rom16_inst_127_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_949 (
  .O(mux_o_949),
  .I0(rom16_inst_143_dout[15]),
  .I1(rom16_inst_159_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_950 (
  .O(mux_o_950),
  .I0(rom16_inst_175_dout[15]),
  .I1(rom16_inst_191_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_951 (
  .O(mux_o_951),
  .I0(rom16_inst_207_dout[15]),
  .I1(rom16_inst_223_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_952 (
  .O(mux_o_952),
  .I0(rom16_inst_239_dout[15]),
  .I1(rom16_inst_255_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_953 (
  .O(mux_o_953),
  .I0(rom16_inst_271_dout[15]),
  .I1(rom16_inst_287_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_954 (
  .O(mux_o_954),
  .I0(rom16_inst_303_dout[15]),
  .I1(rom16_inst_319_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_955 (
  .O(mux_o_955),
  .I0(rom16_inst_335_dout[15]),
  .I1(rom16_inst_351_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_956 (
  .O(mux_o_956),
  .I0(rom16_inst_367_dout[15]),
  .I1(rom16_inst_383_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_957 (
  .O(mux_o_957),
  .I0(rom16_inst_399_dout[15]),
  .I1(rom16_inst_415_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_958 (
  .O(mux_o_958),
  .I0(rom16_inst_431_dout[15]),
  .I1(rom16_inst_447_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_959 (
  .O(mux_o_959),
  .I0(rom16_inst_463_dout[15]),
  .I1(rom16_inst_479_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_960 (
  .O(mux_o_960),
  .I0(rom16_inst_495_dout[15]),
  .I1(rom16_inst_511_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_961 (
  .O(mux_o_961),
  .I0(rom16_inst_527_dout[15]),
  .I1(rom16_inst_543_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_962 (
  .O(mux_o_962),
  .I0(rom16_inst_559_dout[15]),
  .I1(rom16_inst_575_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_963 (
  .O(mux_o_963),
  .I0(rom16_inst_591_dout[15]),
  .I1(rom16_inst_607_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_964 (
  .O(mux_o_964),
  .I0(rom16_inst_623_dout[15]),
  .I1(rom16_inst_639_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_965 (
  .O(mux_o_965),
  .I0(rom16_inst_655_dout[15]),
  .I1(rom16_inst_671_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_966 (
  .O(mux_o_966),
  .I0(rom16_inst_687_dout[15]),
  .I1(rom16_inst_703_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_967 (
  .O(mux_o_967),
  .I0(rom16_inst_719_dout[15]),
  .I1(rom16_inst_735_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_968 (
  .O(mux_o_968),
  .I0(rom16_inst_751_dout[15]),
  .I1(rom16_inst_767_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_969 (
  .O(mux_o_969),
  .I0(rom16_inst_783_dout[15]),
  .I1(rom16_inst_799_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_970 (
  .O(mux_o_970),
  .I0(rom16_inst_815_dout[15]),
  .I1(rom16_inst_831_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_971 (
  .O(mux_o_971),
  .I0(rom16_inst_847_dout[15]),
  .I1(rom16_inst_863_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_972 (
  .O(mux_o_972),
  .I0(rom16_inst_879_dout[15]),
  .I1(rom16_inst_895_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_973 (
  .O(mux_o_973),
  .I0(rom16_inst_911_dout[15]),
  .I1(rom16_inst_927_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_974 (
  .O(mux_o_974),
  .I0(rom16_inst_943_dout[15]),
  .I1(rom16_inst_959_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_975 (
  .O(mux_o_975),
  .I0(rom16_inst_975_dout[15]),
  .I1(rom16_inst_991_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_976 (
  .O(mux_o_976),
  .I0(rom16_inst_1007_dout[15]),
  .I1(rom16_inst_1023_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_977 (
  .O(mux_o_977),
  .I0(mux_o_945),
  .I1(mux_o_946),
  .S0(ad[5])
);
MUX2 mux_inst_978 (
  .O(mux_o_978),
  .I0(mux_o_947),
  .I1(mux_o_948),
  .S0(ad[5])
);
MUX2 mux_inst_979 (
  .O(mux_o_979),
  .I0(mux_o_949),
  .I1(mux_o_950),
  .S0(ad[5])
);
MUX2 mux_inst_980 (
  .O(mux_o_980),
  .I0(mux_o_951),
  .I1(mux_o_952),
  .S0(ad[5])
);
MUX2 mux_inst_981 (
  .O(mux_o_981),
  .I0(mux_o_953),
  .I1(mux_o_954),
  .S0(ad[5])
);
MUX2 mux_inst_982 (
  .O(mux_o_982),
  .I0(mux_o_955),
  .I1(mux_o_956),
  .S0(ad[5])
);
MUX2 mux_inst_983 (
  .O(mux_o_983),
  .I0(mux_o_957),
  .I1(mux_o_958),
  .S0(ad[5])
);
MUX2 mux_inst_984 (
  .O(mux_o_984),
  .I0(mux_o_959),
  .I1(mux_o_960),
  .S0(ad[5])
);
MUX2 mux_inst_985 (
  .O(mux_o_985),
  .I0(mux_o_961),
  .I1(mux_o_962),
  .S0(ad[5])
);
MUX2 mux_inst_986 (
  .O(mux_o_986),
  .I0(mux_o_963),
  .I1(mux_o_964),
  .S0(ad[5])
);
MUX2 mux_inst_987 (
  .O(mux_o_987),
  .I0(mux_o_965),
  .I1(mux_o_966),
  .S0(ad[5])
);
MUX2 mux_inst_988 (
  .O(mux_o_988),
  .I0(mux_o_967),
  .I1(mux_o_968),
  .S0(ad[5])
);
MUX2 mux_inst_989 (
  .O(mux_o_989),
  .I0(mux_o_969),
  .I1(mux_o_970),
  .S0(ad[5])
);
MUX2 mux_inst_990 (
  .O(mux_o_990),
  .I0(mux_o_971),
  .I1(mux_o_972),
  .S0(ad[5])
);
MUX2 mux_inst_991 (
  .O(mux_o_991),
  .I0(mux_o_973),
  .I1(mux_o_974),
  .S0(ad[5])
);
MUX2 mux_inst_992 (
  .O(mux_o_992),
  .I0(mux_o_975),
  .I1(mux_o_976),
  .S0(ad[5])
);
MUX2 mux_inst_993 (
  .O(mux_o_993),
  .I0(mux_o_977),
  .I1(mux_o_978),
  .S0(ad[6])
);
MUX2 mux_inst_994 (
  .O(mux_o_994),
  .I0(mux_o_979),
  .I1(mux_o_980),
  .S0(ad[6])
);
MUX2 mux_inst_995 (
  .O(mux_o_995),
  .I0(mux_o_981),
  .I1(mux_o_982),
  .S0(ad[6])
);
MUX2 mux_inst_996 (
  .O(mux_o_996),
  .I0(mux_o_983),
  .I1(mux_o_984),
  .S0(ad[6])
);
MUX2 mux_inst_997 (
  .O(mux_o_997),
  .I0(mux_o_985),
  .I1(mux_o_986),
  .S0(ad[6])
);
MUX2 mux_inst_998 (
  .O(mux_o_998),
  .I0(mux_o_987),
  .I1(mux_o_988),
  .S0(ad[6])
);
MUX2 mux_inst_999 (
  .O(mux_o_999),
  .I0(mux_o_989),
  .I1(mux_o_990),
  .S0(ad[6])
);
MUX2 mux_inst_1000 (
  .O(mux_o_1000),
  .I0(mux_o_991),
  .I1(mux_o_992),
  .S0(ad[6])
);
MUX2 mux_inst_1001 (
  .O(mux_o_1001),
  .I0(mux_o_993),
  .I1(mux_o_994),
  .S0(ad[7])
);
MUX2 mux_inst_1002 (
  .O(mux_o_1002),
  .I0(mux_o_995),
  .I1(mux_o_996),
  .S0(ad[7])
);
MUX2 mux_inst_1003 (
  .O(mux_o_1003),
  .I0(mux_o_997),
  .I1(mux_o_998),
  .S0(ad[7])
);
MUX2 mux_inst_1004 (
  .O(mux_o_1004),
  .I0(mux_o_999),
  .I1(mux_o_1000),
  .S0(ad[7])
);
MUX2 mux_inst_1005 (
  .O(mux_o_1005),
  .I0(mux_o_1001),
  .I1(mux_o_1002),
  .S0(ad[8])
);
MUX2 mux_inst_1006 (
  .O(mux_o_1006),
  .I0(mux_o_1003),
  .I1(mux_o_1004),
  .S0(ad[8])
);
MUX2 mux_inst_1007 (
  .O(dout[15]),
  .I0(mux_o_1005),
  .I1(mux_o_1006),
  .S0(ad[9])
);
endmodule //inst_mem
